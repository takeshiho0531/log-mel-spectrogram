`timescale	1ns/1ns
module mel_filter_coef # (
    parameter I_BW = 14,
    parameter O_BW = 14
)(
    input clk,
    input rst,
    input [9:0] filter_v, // 0-512
    input signed [I_BW-1:0] data_i, // to adjust timing
    input di_en,
    input is_first_in,
    input is_last_in, // to adjust timing
    output reg signed [O_BW*64-1:0] coef,
    output reg do_en,
    output reg [9:0] out_filter_v,  // 0-512
    output reg signed [O_BW-1:0] data_o,
    output reg is_first_out,
    output reg is_last_out
);
    wire [41:0] non_zero_info_rom [0:512];
    wire [41:0] non_zero_info;

    wire [1:0] non_zero_num;
    wire [5:0] non_zero_idx1;
    wire [5:0] non_zero_idx2;
    wire [9:0] non_zero_data1_addr;
    wire [9:0] non_zero_data2_addr;
    wire signed [15:0] non_zero_data1;
    wire signed [15:0] non_zero_data2;
    reg signed [O_BW*64-1:0] tmp;
    integer i;

    assign non_zero_info = non_zero_info_rom[filter_v];

    assign non_zero_num = non_zero_info[41:40];
    assign non_zero_idx1 = non_zero_info[39:34];
    assign non_zero_idx2 = non_zero_info[33:28];
    assign non_zero_data1_addr = (64-non_zero_idx1)*O_BW;
    assign non_zero_data2_addr = (64-non_zero_idx2)*O_BW;
    assign non_zero_data1 = non_zero_info[27:14];
    assign non_zero_data2 = non_zero_info[13:0];

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            coef <= 0;
            do_en <= 0;
        end else begin
            if (non_zero_num == 0) begin
                do_en <= 0;
                coef <= 0;
                out_filter_v <= filter_v;
                data_o <= data_i;
                do_en<=di_en;
                is_first_out <= is_first_in;
                is_last_out <= is_last_in;
            end
            else if (non_zero_num == 1) begin
                do_en <= 0;
                tmp <= 42'b0;
                for (i=0; i<O_BW; i=i + 1) begin
                    tmp[non_zero_data1_addr-O_BW+i] = non_zero_data1[i];
                end
                coef <= tmp;
                out_filter_v <= filter_v;
                data_o <= data_i;
                do_en<=di_en;
                is_first_out <= is_first_in;
                is_last_out <= is_last_in;
            end
            else if (non_zero_num == 2) begin
                do_en <= 0;
                tmp <= 42'b0;
                for (i=0; i<O_BW; i=i + 1) begin
                    tmp[non_zero_data1_addr-O_BW+i] = non_zero_data1[i];
                    tmp[non_zero_data2_addr-O_BW+i] = non_zero_data2[i];
                end
                coef <= tmp;
                out_filter_v <= filter_v;
                data_o <= data_i;
                do_en <= di_en;
                is_first_out <= is_first_in;
                is_last_out <= is_last_in;
            end
        end    
    end

    assign non_zero_info_rom[0] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[1] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[2] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[3] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[4] = {2'd1, 6'd0, 6'bxxxxxx,14'b00000000001010, 14'bxxxxxxxxxxxxxx}; // 10
    assign non_zero_info_rom[5] = {2'd1, 6'd0, 6'bxxxxxx,14'b00000001001001, 14'bxxxxxxxxxxxxxx}; // 73
    assign non_zero_info_rom[6] = {2'd1, 6'd0, 6'bxxxxxx,14'b00000010001000, 14'bxxxxxxxxxxxxxx}; // 136
    assign non_zero_info_rom[7] = {2'd2, 6'd0, 6'd1,14'b00000010100100, 14'b00000000010001}; // 164, 17
    assign non_zero_info_rom[8] = {2'd2, 6'd0, 6'd1,14'b00000001100110, 14'b00000001010000}; // 102, 80
    assign non_zero_info_rom[9] = {2'd2, 6'd0, 6'd1,14'b00000000100111, 14'b00000010001111}; // 39, 143
    assign non_zero_info_rom[10] = {2'd2, 6'd1, 6'd2,14'b00000010011101, 14'b00000000011000}; // 157, 24
    assign non_zero_info_rom[11] = {2'd2, 6'd1, 6'd2,14'b00000001011110, 14'b00000001010111}; // 94, 87
    assign non_zero_info_rom[12] = {2'd2, 6'd1, 6'd2,14'b00000000011111, 14'b00000010010110}; // 31, 150
    assign non_zero_info_rom[13] = {2'd2, 6'd2, 6'd3,14'b00000010010110, 14'b00000000011111}; // 150, 31
    assign non_zero_info_rom[14] = {2'd2, 6'd2, 6'd3,14'b00000001010111, 14'b00000001011110}; // 87, 94
    assign non_zero_info_rom[15] = {2'd2, 6'd2, 6'd3,14'b00000000011000, 14'b00000010011101}; // 24, 157
    assign non_zero_info_rom[16] = {2'd2, 6'd3, 6'd4,14'b00000010001111, 14'b00000000100111}; // 143, 39
    assign non_zero_info_rom[17] = {2'd2, 6'd3, 6'd4,14'b00000001010000, 14'b00000001100101}; // 80, 101
    assign non_zero_info_rom[18] = {2'd2, 6'd3, 6'd4,14'b00000000010001, 14'b00000010100100}; // 17, 164
    assign non_zero_info_rom[19] = {2'd2, 6'd4, 6'd5,14'b00000010001000, 14'b00000000101110}; // 136, 46
    assign non_zero_info_rom[20] = {2'd2, 6'd4, 6'd5,14'b00000001001001, 14'b00000001101101}; // 73, 109
    assign non_zero_info_rom[21] = {2'd2, 6'd4, 6'd5,14'b00000000001010, 14'b00000010101100}; // 10, 172
    assign non_zero_info_rom[22] = {2'd2, 6'd5, 6'd6,14'b00000010000001, 14'b00000000110101}; // 129, 53
    assign non_zero_info_rom[23] = {2'd2, 6'd5, 6'd6,14'b00000001000010, 14'b00000001110100}; // 66, 116
    assign non_zero_info_rom[24] = {2'd2, 6'd5, 6'd6,14'b00000000000011, 14'b00000010110011}; // 3, 179
    assign non_zero_info_rom[25] = {2'd2, 6'd6, 6'd7,14'b00000001111010, 14'b00000000111100}; // 122, 60
    assign non_zero_info_rom[26] = {2'd2, 6'd6, 6'd7,14'b00000000111011, 14'b00000001111011}; // 59, 123
    assign non_zero_info_rom[27] = {2'd2, 6'd7, 6'd8,14'b00000010110001, 14'b00000000000100}; // 177, 4
    assign non_zero_info_rom[28] = {2'd2, 6'd7, 6'd8,14'b00000001110011, 14'b00000001000011}; // 115, 67
    assign non_zero_info_rom[29] = {2'd2, 6'd7, 6'd8,14'b00000000110100, 14'b00000010000010}; // 52, 130
    assign non_zero_info_rom[30] = {2'd2, 6'd8, 6'd9,14'b00000010101010, 14'b00000000001011}; // 170, 11
    assign non_zero_info_rom[31] = {2'd2, 6'd8, 6'd9,14'b00000001101011, 14'b00000001001010}; // 107, 74
    assign non_zero_info_rom[32] = {2'd2, 6'd8, 6'd9,14'b00000000101100, 14'b00000010001001}; // 44, 137
    assign non_zero_info_rom[33] = {2'd2, 6'd9, 6'd10,14'b00000010100011, 14'b00000000010010}; // 163, 18
    assign non_zero_info_rom[34] = {2'd2, 6'd9, 6'd10,14'b00000001100100, 14'b00000001010001}; // 100, 81
    assign non_zero_info_rom[35] = {2'd2, 6'd9, 6'd10,14'b00000000100101, 14'b00000010010000}; // 37, 144
    assign non_zero_info_rom[36] = {2'd2, 6'd10, 6'd11,14'b00000010011100, 14'b00000000011010}; // 156, 26
    assign non_zero_info_rom[37] = {2'd2, 6'd10, 6'd11,14'b00000001011101, 14'b00000001011000}; // 93, 88
    assign non_zero_info_rom[38] = {2'd2, 6'd10, 6'd11,14'b00000000011110, 14'b00000010010111}; // 30, 151
    assign non_zero_info_rom[39] = {2'd2, 6'd11, 6'd12,14'b00000010010101, 14'b00000000100001}; // 149, 33
    assign non_zero_info_rom[40] = {2'd2, 6'd11, 6'd12,14'b00000001010110, 14'b00000001100000}; // 86, 96
    assign non_zero_info_rom[41] = {2'd2, 6'd11, 6'd12,14'b00000000010111, 14'b00000010011111}; // 23, 159
    assign non_zero_info_rom[42] = {2'd2, 6'd12, 6'd13,14'b00000010001110, 14'b00000000101000}; // 142, 40
    assign non_zero_info_rom[43] = {2'd2, 6'd12, 6'd13,14'b00000001001111, 14'b00000001100111}; // 79, 103
    assign non_zero_info_rom[44] = {2'd2, 6'd12, 6'd13,14'b00000000010000, 14'b00000010100110}; // 16, 166
    assign non_zero_info_rom[45] = {2'd2, 6'd13, 6'd14,14'b00000010000111, 14'b00000000101111}; // 135, 47
    assign non_zero_info_rom[46] = {2'd2, 6'd13, 6'd14,14'b00000001001000, 14'b00000001101110}; // 72, 110
    assign non_zero_info_rom[47] = {2'd2, 6'd13, 6'd14,14'b00000000001001, 14'b00000010101101}; // 9, 173
    assign non_zero_info_rom[48] = {2'd2, 6'd14, 6'd15,14'b00000010000000, 14'b00000000110110}; // 128, 54
    assign non_zero_info_rom[49] = {2'd2, 6'd14, 6'd15,14'b00000001000001, 14'b00000001110101}; // 65, 117
    assign non_zero_info_rom[50] = {2'd2, 6'd14, 6'd15,14'b00000000000010, 14'b00000010110100}; // 2, 180
    assign non_zero_info_rom[51] = {2'd2, 6'd15, 6'd16,14'b00000001111000, 14'b00000000111101}; // 120, 61
    assign non_zero_info_rom[52] = {2'd2, 6'd15, 6'd16,14'b00000000111010, 14'b00000001111100}; // 58, 124
    assign non_zero_info_rom[53] = {2'd2, 6'd16, 6'd17,14'b00000010110000, 14'b00000000000101}; // 176, 5
    assign non_zero_info_rom[54] = {2'd2, 6'd16, 6'd17,14'b00000001110001, 14'b00000001000100}; // 113, 68
    assign non_zero_info_rom[55] = {2'd2, 6'd16, 6'd17,14'b00000000110010, 14'b00000010000011}; // 50, 131
    assign non_zero_info_rom[56] = {2'd2, 6'd17, 6'd18,14'b00000010101001, 14'b00000000001101}; // 169, 13
    assign non_zero_info_rom[57] = {2'd2, 6'd17, 6'd18,14'b00000001101010, 14'b00000001001011}; // 106, 75
    assign non_zero_info_rom[58] = {2'd2, 6'd17, 6'd18,14'b00000000101011, 14'b00000010001010}; // 43, 138
    assign non_zero_info_rom[59] = {2'd2, 6'd18, 6'd19,14'b00000010100010, 14'b00000000010100}; // 162, 20
    assign non_zero_info_rom[60] = {2'd2, 6'd18, 6'd19,14'b00000001100011, 14'b00000001010010}; // 99, 82
    assign non_zero_info_rom[61] = {2'd2, 6'd18, 6'd19,14'b00000000100100, 14'b00000010010001}; // 36, 145
    assign non_zero_info_rom[62] = {2'd2, 6'd19, 6'd20,14'b00000010011011, 14'b00000000011010}; // 155, 26
    assign non_zero_info_rom[63] = {2'd2, 6'd19, 6'd20,14'b00000001011100, 14'b00000001010110}; // 92, 86
    assign non_zero_info_rom[64] = {2'd2, 6'd19, 6'd20,14'b00000000011110, 14'b00000010010011}; // 30, 147
    assign non_zero_info_rom[65] = {2'd2, 6'd20, 6'd21,14'b00000010010010, 14'b00000000011100}; // 146, 28
    assign non_zero_info_rom[66] = {2'd2, 6'd20, 6'd21,14'b00000001011000, 14'b00000001010011}; // 88, 83
    assign non_zero_info_rom[67] = {2'd2, 6'd20, 6'd21,14'b00000000011111, 14'b00000010001001}; // 31, 137
    assign non_zero_info_rom[68] = {2'd2, 6'd21, 6'd22,14'b00000010001111, 14'b00000000010110}; // 143, 22
    assign non_zero_info_rom[69] = {2'd2, 6'd21, 6'd22,14'b00000001011011, 14'b00000001001000}; // 91, 72
    assign non_zero_info_rom[70] = {2'd2, 6'd21, 6'd22,14'b00000000101000, 14'b00000001111001}; // 40, 121
    assign non_zero_info_rom[71] = {2'd2, 6'd22, 6'd23,14'b00000010010100, 14'b00000000001011}; // 148, 11
    assign non_zero_info_rom[72] = {2'd2, 6'd22, 6'd23,14'b00000001100101, 14'b00000000111000}; // 101, 56
    assign non_zero_info_rom[73] = {2'd2, 6'd22, 6'd23,14'b00000000110110, 14'b00000001100101}; // 54, 101
    assign non_zero_info_rom[74] = {2'd2, 6'd22, 6'd23,14'b00000000000110, 14'b00000010010010}; // 6, 146
    assign non_zero_info_rom[75] = {2'd2, 6'd23, 6'd24,14'b00000001110011, 14'b00000000100100}; // 115, 36
    assign non_zero_info_rom[76] = {2'd2, 6'd23, 6'd24,14'b00000001001000, 14'b00000001001101}; // 72, 77
    assign non_zero_info_rom[77] = {2'd2, 6'd23, 6'd24,14'b00000000011101, 14'b00000001110110}; // 29, 118
    assign non_zero_info_rom[78] = {2'd2, 6'd24, 6'd25,14'b00000010000100, 14'b00000000001101}; // 132, 13
    assign non_zero_info_rom[79] = {2'd2, 6'd24, 6'd25,14'b00000001011101, 14'b00000000110010}; // 93, 50
    assign non_zero_info_rom[80] = {2'd2, 6'd24, 6'd25,14'b00000000110101, 14'b00000001011000}; // 53, 88
    assign non_zero_info_rom[81] = {2'd2, 6'd24, 6'd25,14'b00000000001110, 14'b00000001111101}; // 14, 125
    assign non_zero_info_rom[82] = {2'd2, 6'd25, 6'd26,14'b00000001110100, 14'b00000000010110}; // 116, 22
    assign non_zero_info_rom[83] = {2'd2, 6'd25, 6'd26,14'b00000001010000, 14'b00000000111000}; // 80, 56
    assign non_zero_info_rom[84] = {2'd2, 6'd25, 6'd26,14'b00000000101100, 14'b00000001011010}; // 44, 90
    assign non_zero_info_rom[85] = {2'd2, 6'd25, 6'd26,14'b00000000001000, 14'b00000001111100}; // 8, 124
    assign non_zero_info_rom[86] = {2'd2, 6'd26, 6'd27,14'b00000001101011, 14'b00000000011000}; // 107, 24
    assign non_zero_info_rom[87] = {2'd2, 6'd26, 6'd27,14'b00000001001011, 14'b00000000110111}; // 75, 55
    assign non_zero_info_rom[88] = {2'd2, 6'd26, 6'd27,14'b00000000101010, 14'b00000001010110}; // 42, 86
    assign non_zero_info_rom[89] = {2'd2, 6'd26, 6'd27,14'b00000000001010, 14'b00000001110101}; // 10, 117
    assign non_zero_info_rom[90] = {2'd2, 6'd27, 6'd28,14'b00000001101001, 14'b00000000010100}; // 105, 20
    assign non_zero_info_rom[91] = {2'd2, 6'd27, 6'd28,14'b00000001001100, 14'b00000000110000}; // 76, 48
    assign non_zero_info_rom[92] = {2'd2, 6'd27, 6'd28,14'b00000000101110, 14'b00000001001101}; // 46, 77
    assign non_zero_info_rom[93] = {2'd2, 6'd27, 6'd28,14'b00000000010000, 14'b00000001101001}; // 16, 105
    assign non_zero_info_rom[94] = {2'd2, 6'd28, 6'd29,14'b00000001101100, 14'b00000000001100}; // 108, 12
    assign non_zero_info_rom[95] = {2'd2, 6'd28, 6'd29,14'b00000001010001, 14'b00000000100110}; // 81, 38
    assign non_zero_info_rom[96] = {2'd2, 6'd28, 6'd29,14'b00000000110110, 14'b00000000111111}; // 54, 63
    assign non_zero_info_rom[97] = {2'd2, 6'd28, 6'd29,14'b00000000011011, 14'b00000001011001}; // 27, 89
    assign non_zero_info_rom[98] = {2'd2, 6'd29, 6'd30,14'b00000001110011, 14'b00000000000000}; // 115, 0
    assign non_zero_info_rom[99] = {2'd2, 6'd29, 6'd30,14'b00000001011010, 14'b00000000011000}; // 90, 24
    assign non_zero_info_rom[100] = {2'd2, 6'd29, 6'd30,14'b00000001000010, 14'b00000000101111}; // 66, 47
    assign non_zero_info_rom[101] = {2'd2, 6'd29, 6'd30,14'b00000000101001, 14'b00000001000111}; // 41, 71
    assign non_zero_info_rom[102] = {2'd2, 6'd29, 6'd30,14'b00000000010000, 14'b00000001011110}; // 16, 94
    assign non_zero_info_rom[103] = {2'd2, 6'd30, 6'd31,14'b00000001100110, 14'b00000000000111}; // 102, 7
    assign non_zero_info_rom[104] = {2'd2, 6'd30, 6'd31,14'b00000001010000, 14'b00000000011101}; // 80, 29
    assign non_zero_info_rom[105] = {2'd2, 6'd30, 6'd31,14'b00000000111001, 14'b00000000110010}; // 57, 50
    assign non_zero_info_rom[106] = {2'd2, 6'd30, 6'd31,14'b00000000100011, 14'b00000001000111}; // 35, 71
    assign non_zero_info_rom[107] = {2'd2, 6'd30, 6'd31,14'b00000000001100, 14'b00000001011101}; // 12, 93
    assign non_zero_info_rom[108] = {2'd2, 6'd31, 6'd32,14'b00000001100000, 14'b00000000001001}; // 96, 9
    assign non_zero_info_rom[109] = {2'd2, 6'd31, 6'd32,14'b00000001001011, 14'b00000000011100}; // 75, 28
    assign non_zero_info_rom[110] = {2'd2, 6'd31, 6'd32,14'b00000000110111, 14'b00000000110000}; // 55, 48
    assign non_zero_info_rom[111] = {2'd2, 6'd31, 6'd32,14'b00000000100010, 14'b00000001000011}; // 34, 67
    assign non_zero_info_rom[112] = {2'd2, 6'd31, 6'd32,14'b00000000001110, 14'b00000001010111}; // 14, 87
    assign non_zero_info_rom[113] = {2'd2, 6'd32, 6'd33,14'b00000001011110, 14'b00000000000110}; // 94, 6
    assign non_zero_info_rom[114] = {2'd2, 6'd32, 6'd33,14'b00000001001011, 14'b00000000011000}; // 75, 24
    assign non_zero_info_rom[115] = {2'd2, 6'd32, 6'd33,14'b00000000111001, 14'b00000000101001}; // 57, 41
    assign non_zero_info_rom[116] = {2'd2, 6'd32, 6'd33,14'b00000000100110, 14'b00000000111011}; // 38, 59
    assign non_zero_info_rom[117] = {2'd2, 6'd32, 6'd33,14'b00000000010011, 14'b00000001001101}; // 19, 77
    assign non_zero_info_rom[118] = {2'd2, 6'd32, 6'd33,14'b00000000000001, 14'b00000001011111}; // 1, 95
    assign non_zero_info_rom[119] = {2'd2, 6'd33, 6'd34,14'b00000001001111, 14'b00000000010000}; // 79, 16
    assign non_zero_info_rom[120] = {2'd2, 6'd33, 6'd34,14'b00000000111110, 14'b00000000100000}; // 62, 32
    assign non_zero_info_rom[121] = {2'd2, 6'd33, 6'd34,14'b00000000101101, 14'b00000000110000}; // 45, 48
    assign non_zero_info_rom[122] = {2'd2, 6'd33, 6'd34,14'b00000000011100, 14'b00000001000000}; // 28, 64
    assign non_zero_info_rom[123] = {2'd2, 6'd33, 6'd34,14'b00000000001011, 14'b00000001010000}; // 11, 80
    assign non_zero_info_rom[124] = {2'd2, 6'd34, 6'd35,14'b00000001010110, 14'b00000000000101}; // 86, 5
    assign non_zero_info_rom[125] = {2'd2, 6'd34, 6'd35,14'b00000001000110, 14'b00000000010100}; // 70, 20
    assign non_zero_info_rom[126] = {2'd2, 6'd34, 6'd35,14'b00000000110111, 14'b00000000100011}; // 55, 35
    assign non_zero_info_rom[127] = {2'd2, 6'd34, 6'd35,14'b00000000100111, 14'b00000000110001}; // 39, 49
    assign non_zero_info_rom[128] = {2'd2, 6'd34, 6'd35,14'b00000000011000, 14'b00000001000000}; // 24, 64
    assign non_zero_info_rom[129] = {2'd2, 6'd34, 6'd35,14'b00000000001000, 14'b00000001001111}; // 8, 79
    assign non_zero_info_rom[130] = {2'd2, 6'd35, 6'd36,14'b00000001010001, 14'b00000000000110}; // 81, 6
    assign non_zero_info_rom[131] = {2'd2, 6'd35, 6'd36,14'b00000001000010, 14'b00000000010100}; // 66, 20
    assign non_zero_info_rom[132] = {2'd2, 6'd35, 6'd36,14'b00000000110100, 14'b00000000100001}; // 52, 33
    assign non_zero_info_rom[133] = {2'd2, 6'd35, 6'd36,14'b00000000100110, 14'b00000000101110}; // 38, 46
    assign non_zero_info_rom[134] = {2'd2, 6'd35, 6'd36,14'b00000000011000, 14'b00000000111100}; // 24, 60
    assign non_zero_info_rom[135] = {2'd2, 6'd35, 6'd36,14'b00000000001010, 14'b00000001001001}; // 10, 73
    assign non_zero_info_rom[136] = {2'd2, 6'd36, 6'd37,14'b00000001001111, 14'b00000000000011}; // 79, 3
    assign non_zero_info_rom[137] = {2'd2, 6'd36, 6'd37,14'b00000001000011, 14'b00000000010000}; // 67, 16
    assign non_zero_info_rom[138] = {2'd2, 6'd36, 6'd37,14'b00000000110110, 14'b00000000011100}; // 54, 28
    assign non_zero_info_rom[139] = {2'd2, 6'd36, 6'd37,14'b00000000101001, 14'b00000000101000}; // 41, 40
    assign non_zero_info_rom[140] = {2'd2, 6'd36, 6'd37,14'b00000000011100, 14'b00000000110101}; // 28, 53
    assign non_zero_info_rom[141] = {2'd2, 6'd36, 6'd37,14'b00000000001111, 14'b00000001000001}; // 15, 65
    assign non_zero_info_rom[142] = {2'd2, 6'd36, 6'd37,14'b00000000000010, 14'b00000001001101}; // 2, 77
    assign non_zero_info_rom[143] = {2'd2, 6'd37, 6'd38,14'b00000001000110, 14'b00000000001001}; // 70, 9
    assign non_zero_info_rom[144] = {2'd2, 6'd37, 6'd38,14'b00000000111010, 14'b00000000010100}; // 58, 20
    assign non_zero_info_rom[145] = {2'd2, 6'd37, 6'd38,14'b00000000101110, 14'b00000000100000}; // 46, 32
    assign non_zero_info_rom[146] = {2'd2, 6'd37, 6'd38,14'b00000000100011, 14'b00000000101011}; // 35, 43
    assign non_zero_info_rom[147] = {2'd2, 6'd37, 6'd38,14'b00000000010111, 14'b00000000110110}; // 23, 54
    assign non_zero_info_rom[148] = {2'd2, 6'd37, 6'd38,14'b00000000001011, 14'b00000001000001}; // 11, 65
    assign non_zero_info_rom[149] = {2'd2, 6'd38, 6'd39,14'b00000001001011, 14'b00000000000001}; // 75, 1
    assign non_zero_info_rom[150] = {2'd2, 6'd38, 6'd39,14'b00000001000000, 14'b00000000001011}; // 64, 11
    assign non_zero_info_rom[151] = {2'd2, 6'd38, 6'd39,14'b00000000110110, 14'b00000000010101}; // 54, 21
    assign non_zero_info_rom[152] = {2'd2, 6'd38, 6'd39,14'b00000000101011, 14'b00000000011111}; // 43, 31
    assign non_zero_info_rom[153] = {2'd2, 6'd38, 6'd39,14'b00000000100000, 14'b00000000101001}; // 32, 41
    assign non_zero_info_rom[154] = {2'd2, 6'd38, 6'd39,14'b00000000010110, 14'b00000000110011}; // 22, 51
    assign non_zero_info_rom[155] = {2'd2, 6'd38, 6'd39,14'b00000000001011, 14'b00000000111110}; // 11, 62
    assign non_zero_info_rom[156] = {2'd2, 6'd38, 6'd39,14'b00000000000000, 14'b00000001001000}; // 0, 72
    assign non_zero_info_rom[157] = {2'd2, 6'd39, 6'd40,14'b00000000111111, 14'b00000000001001}; // 63, 9
    assign non_zero_info_rom[158] = {2'd2, 6'd39, 6'd40,14'b00000000110101, 14'b00000000010010}; // 53, 18
    assign non_zero_info_rom[159] = {2'd2, 6'd39, 6'd40,14'b00000000101011, 14'b00000000011011}; // 43, 27
    assign non_zero_info_rom[160] = {2'd2, 6'd39, 6'd40,14'b00000000100010, 14'b00000000100101}; // 34, 37
    assign non_zero_info_rom[161] = {2'd2, 6'd39, 6'd40,14'b00000000011000, 14'b00000000101110}; // 24, 46
    assign non_zero_info_rom[162] = {2'd2, 6'd39, 6'd40,14'b00000000001110, 14'b00000000110111}; // 14, 55
    assign non_zero_info_rom[163] = {2'd2, 6'd39, 6'd40,14'b00000000000101, 14'b00000001000001}; // 5, 65
    assign non_zero_info_rom[164] = {2'd2, 6'd40, 6'd41,14'b00000001000000, 14'b00000000000100}; // 64, 4
    assign non_zero_info_rom[165] = {2'd2, 6'd40, 6'd41,14'b00000000110111, 14'b00000000001101}; // 55, 13
    assign non_zero_info_rom[166] = {2'd2, 6'd40, 6'd41,14'b00000000101111, 14'b00000000010101}; // 47, 21
    assign non_zero_info_rom[167] = {2'd2, 6'd40, 6'd41,14'b00000000100110, 14'b00000000011110}; // 38, 30
    assign non_zero_info_rom[168] = {2'd2, 6'd40, 6'd41,14'b00000000011101, 14'b00000000100110}; // 29, 38
    assign non_zero_info_rom[169] = {2'd2, 6'd40, 6'd41,14'b00000000010100, 14'b00000000101111}; // 20, 47
    assign non_zero_info_rom[170] = {2'd2, 6'd40, 6'd41,14'b00000000001011, 14'b00000000110111}; // 11, 55
    assign non_zero_info_rom[171] = {2'd2, 6'd40, 6'd41,14'b00000000000010, 14'b00000001000000}; // 2, 64
    assign non_zero_info_rom[172] = {2'd2, 6'd41, 6'd42,14'b00000000111100, 14'b00000000000110}; // 60, 6
    assign non_zero_info_rom[173] = {2'd2, 6'd41, 6'd42,14'b00000000110100, 14'b00000000001101}; // 52, 13
    assign non_zero_info_rom[174] = {2'd2, 6'd41, 6'd42,14'b00000000101100, 14'b00000000010101}; // 44, 21
    assign non_zero_info_rom[175] = {2'd2, 6'd41, 6'd42,14'b00000000100100, 14'b00000000011101}; // 36, 29
    assign non_zero_info_rom[176] = {2'd2, 6'd41, 6'd42,14'b00000000011011, 14'b00000000100101}; // 27, 37
    assign non_zero_info_rom[177] = {2'd2, 6'd41, 6'd42,14'b00000000010011, 14'b00000000101100}; // 19, 44
    assign non_zero_info_rom[178] = {2'd2, 6'd41, 6'd42,14'b00000000001011, 14'b00000000110100}; // 11, 52
    assign non_zero_info_rom[179] = {2'd2, 6'd41, 6'd42,14'b00000000000011, 14'b00000000111100}; // 3, 60
    assign non_zero_info_rom[180] = {2'd2, 6'd42, 6'd43,14'b00000000111010, 14'b00000000000100}; // 58, 4
    assign non_zero_info_rom[181] = {2'd2, 6'd42, 6'd43,14'b00000000110011, 14'b00000000001011}; // 51, 11
    assign non_zero_info_rom[182] = {2'd2, 6'd42, 6'd43,14'b00000000101100, 14'b00000000010010}; // 44, 18
    assign non_zero_info_rom[183] = {2'd2, 6'd42, 6'd43,14'b00000000100100, 14'b00000000011001}; // 36, 25
    assign non_zero_info_rom[184] = {2'd2, 6'd42, 6'd43,14'b00000000011101, 14'b00000000100000}; // 29, 32
    assign non_zero_info_rom[185] = {2'd2, 6'd42, 6'd43,14'b00000000010110, 14'b00000000100111}; // 22, 39
    assign non_zero_info_rom[186] = {2'd2, 6'd42, 6'd43,14'b00000000001110, 14'b00000000101110}; // 14, 46
    assign non_zero_info_rom[187] = {2'd2, 6'd42, 6'd43,14'b00000000000111, 14'b00000000110101}; // 7, 53
    assign non_zero_info_rom[188] = {2'd2, 6'd43, 6'd44,14'b00000000111100, 14'b00000000000000}; // 60, 0
    assign non_zero_info_rom[189] = {2'd2, 6'd43, 6'd44,14'b00000000110101, 14'b00000000000111}; // 53, 7
    assign non_zero_info_rom[190] = {2'd2, 6'd43, 6'd44,14'b00000000101110, 14'b00000000001101}; // 46, 13
    assign non_zero_info_rom[191] = {2'd2, 6'd43, 6'd44,14'b00000000101000, 14'b00000000010100}; // 40, 20
    assign non_zero_info_rom[192] = {2'd2, 6'd43, 6'd44,14'b00000000100001, 14'b00000000011010}; // 33, 26
    assign non_zero_info_rom[193] = {2'd2, 6'd43, 6'd44,14'b00000000011010, 14'b00000000100000}; // 26, 32
    assign non_zero_info_rom[194] = {2'd2, 6'd43, 6'd44,14'b00000000010011, 14'b00000000100111}; // 19, 39
    assign non_zero_info_rom[195] = {2'd2, 6'd43, 6'd44,14'b00000000001101, 14'b00000000101101}; // 13, 45
    assign non_zero_info_rom[196] = {2'd2, 6'd43, 6'd44,14'b00000000000110, 14'b00000000110011}; // 6, 51
    assign non_zero_info_rom[197] = {2'd2, 6'd44, 6'd45,14'b00000000111001, 14'b00000000000001}; // 57, 1
    assign non_zero_info_rom[198] = {2'd2, 6'd44, 6'd45,14'b00000000110011, 14'b00000000000110}; // 51, 6
    assign non_zero_info_rom[199] = {2'd2, 6'd44, 6'd45,14'b00000000101100, 14'b00000000001100}; // 44, 12
    assign non_zero_info_rom[200] = {2'd2, 6'd44, 6'd45,14'b00000000100110, 14'b00000000010010}; // 38, 18
    assign non_zero_info_rom[201] = {2'd2, 6'd44, 6'd45,14'b00000000100000, 14'b00000000011000}; // 32, 24
    assign non_zero_info_rom[202] = {2'd2, 6'd44, 6'd45,14'b00000000011010, 14'b00000000011110}; // 26, 30
    assign non_zero_info_rom[203] = {2'd2, 6'd44, 6'd45,14'b00000000010100, 14'b00000000100100}; // 20, 36
    assign non_zero_info_rom[204] = {2'd2, 6'd44, 6'd45,14'b00000000001110, 14'b00000000101001}; // 14, 41
    assign non_zero_info_rom[205] = {2'd2, 6'd44, 6'd45,14'b00000000001000, 14'b00000000101111}; // 8, 47
    assign non_zero_info_rom[206] = {2'd2, 6'd44, 6'd45,14'b00000000000010, 14'b00000000110101}; // 2, 53
    assign non_zero_info_rom[207] = {2'd2, 6'd45, 6'd46,14'b00000000110011, 14'b00000000000100}; // 51, 4
    assign non_zero_info_rom[208] = {2'd2, 6'd45, 6'd46,14'b00000000101101, 14'b00000000001001}; // 45, 9
    assign non_zero_info_rom[209] = {2'd2, 6'd45, 6'd46,14'b00000000100111, 14'b00000000001110}; // 39, 14
    assign non_zero_info_rom[210] = {2'd2, 6'd45, 6'd46,14'b00000000100010, 14'b00000000010100}; // 34, 20
    assign non_zero_info_rom[211] = {2'd2, 6'd45, 6'd46,14'b00000000011100, 14'b00000000011001}; // 28, 25
    assign non_zero_info_rom[212] = {2'd2, 6'd45, 6'd46,14'b00000000010111, 14'b00000000011110}; // 23, 30
    assign non_zero_info_rom[213] = {2'd2, 6'd45, 6'd46,14'b00000000010001, 14'b00000000100100}; // 17, 36
    assign non_zero_info_rom[214] = {2'd2, 6'd45, 6'd46,14'b00000000001100, 14'b00000000101001}; // 12, 41
    assign non_zero_info_rom[215] = {2'd2, 6'd45, 6'd46,14'b00000000000110, 14'b00000000101110}; // 6, 46
    assign non_zero_info_rom[216] = {2'd2, 6'd45, 6'd46,14'b00000000000001, 14'b00000000110100}; // 1, 52
    assign non_zero_info_rom[217] = {2'd2, 6'd46, 6'd47,14'b00000000110000, 14'b00000000000100}; // 48, 4
    assign non_zero_info_rom[218] = {2'd2, 6'd46, 6'd47,14'b00000000101010, 14'b00000000001001}; // 42, 9
    assign non_zero_info_rom[219] = {2'd2, 6'd46, 6'd47,14'b00000000100101, 14'b00000000001110}; // 37, 14
    assign non_zero_info_rom[220] = {2'd2, 6'd46, 6'd47,14'b00000000100000, 14'b00000000010011}; // 32, 19
    assign non_zero_info_rom[221] = {2'd2, 6'd46, 6'd47,14'b00000000011011, 14'b00000000011000}; // 27, 24
    assign non_zero_info_rom[222] = {2'd2, 6'd46, 6'd47,14'b00000000010110, 14'b00000000011101}; // 22, 29
    assign non_zero_info_rom[223] = {2'd2, 6'd46, 6'd47,14'b00000000010001, 14'b00000000100001}; // 17, 33
    assign non_zero_info_rom[224] = {2'd2, 6'd46, 6'd47,14'b00000000001100, 14'b00000000100110}; // 12, 38
    assign non_zero_info_rom[225] = {2'd2, 6'd46, 6'd47,14'b00000000000111, 14'b00000000101011}; // 7, 43
    assign non_zero_info_rom[226] = {2'd2, 6'd46, 6'd47,14'b00000000000010, 14'b00000000110000}; // 2, 48
    assign non_zero_info_rom[227] = {2'd2, 6'd47, 6'd48,14'b00000000101111, 14'b00000000000011}; // 47, 3
    assign non_zero_info_rom[228] = {2'd2, 6'd47, 6'd48,14'b00000000101010, 14'b00000000000111}; // 42, 7
    assign non_zero_info_rom[229] = {2'd2, 6'd47, 6'd48,14'b00000000100110, 14'b00000000001100}; // 38, 12
    assign non_zero_info_rom[230] = {2'd2, 6'd47, 6'd48,14'b00000000100001, 14'b00000000010000}; // 33, 16
    assign non_zero_info_rom[231] = {2'd2, 6'd47, 6'd48,14'b00000000011100, 14'b00000000010100}; // 28, 20
    assign non_zero_info_rom[232] = {2'd2, 6'd47, 6'd48,14'b00000000011000, 14'b00000000011001}; // 24, 25
    assign non_zero_info_rom[233] = {2'd2, 6'd47, 6'd48,14'b00000000010011, 14'b00000000011101}; // 19, 29
    assign non_zero_info_rom[234] = {2'd2, 6'd47, 6'd48,14'b00000000001111, 14'b00000000100010}; // 15, 34
    assign non_zero_info_rom[235] = {2'd2, 6'd47, 6'd48,14'b00000000001010, 14'b00000000100110}; // 10, 38
    assign non_zero_info_rom[236] = {2'd2, 6'd47, 6'd48,14'b00000000000101, 14'b00000000101010}; // 5, 42
    assign non_zero_info_rom[237] = {2'd2, 6'd47, 6'd48,14'b00000000000001, 14'b00000000101111}; // 1, 47
    assign non_zero_info_rom[238] = {2'd2, 6'd48, 6'd49,14'b00000000101100, 14'b00000000000011}; // 44, 3
    assign non_zero_info_rom[239] = {2'd2, 6'd48, 6'd49,14'b00000000101000, 14'b00000000000111}; // 40, 7
    assign non_zero_info_rom[240] = {2'd2, 6'd48, 6'd49,14'b00000000100100, 14'b00000000001011}; // 36, 11
    assign non_zero_info_rom[241] = {2'd2, 6'd48, 6'd49,14'b00000000011111, 14'b00000000001111}; // 31, 15
    assign non_zero_info_rom[242] = {2'd2, 6'd48, 6'd49,14'b00000000011011, 14'b00000000010011}; // 27, 19
    assign non_zero_info_rom[243] = {2'd2, 6'd48, 6'd49,14'b00000000010111, 14'b00000000010111}; // 23, 23
    assign non_zero_info_rom[244] = {2'd2, 6'd48, 6'd49,14'b00000000010011, 14'b00000000011011}; // 19, 27
    assign non_zero_info_rom[245] = {2'd2, 6'd48, 6'd49,14'b00000000001111, 14'b00000000011111}; // 15, 31
    assign non_zero_info_rom[246] = {2'd2, 6'd48, 6'd49,14'b00000000001010, 14'b00000000100011}; // 10, 35
    assign non_zero_info_rom[247] = {2'd2, 6'd48, 6'd49,14'b00000000000110, 14'b00000000100111}; // 6, 39
    assign non_zero_info_rom[248] = {2'd2, 6'd48, 6'd49,14'b00000000000010, 14'b00000000101100}; // 2, 44
    assign non_zero_info_rom[249] = {2'd2, 6'd49, 6'd50,14'b00000000101011, 14'b00000000000010}; // 43, 2
    assign non_zero_info_rom[250] = {2'd2, 6'd49, 6'd50,14'b00000000100111, 14'b00000000000110}; // 39, 6
    assign non_zero_info_rom[251] = {2'd2, 6'd49, 6'd50,14'b00000000100100, 14'b00000000001001}; // 36, 9
    assign non_zero_info_rom[252] = {2'd2, 6'd49, 6'd50,14'b00000000100000, 14'b00000000001101}; // 32, 13
    assign non_zero_info_rom[253] = {2'd2, 6'd49, 6'd50,14'b00000000011100, 14'b00000000010001}; // 28, 17
    assign non_zero_info_rom[254] = {2'd2, 6'd49, 6'd50,14'b00000000011000, 14'b00000000010100}; // 24, 20
    assign non_zero_info_rom[255] = {2'd2, 6'd49, 6'd50,14'b00000000010100, 14'b00000000011000}; // 20, 24
    assign non_zero_info_rom[256] = {2'd2, 6'd49, 6'd50,14'b00000000010000, 14'b00000000011100}; // 16, 28
    assign non_zero_info_rom[257] = {2'd2, 6'd49, 6'd50,14'b00000000001101, 14'b00000000011111}; // 13, 31
    assign non_zero_info_rom[258] = {2'd2, 6'd49, 6'd50,14'b00000000001001, 14'b00000000100011}; // 9, 35
    assign non_zero_info_rom[259] = {2'd2, 6'd49, 6'd50,14'b00000000000101, 14'b00000000100111}; // 5, 39
    assign non_zero_info_rom[260] = {2'd2, 6'd49, 6'd50,14'b00000000000001, 14'b00000000101010}; // 1, 42
    assign non_zero_info_rom[261] = {2'd2, 6'd50, 6'd51,14'b00000000101001, 14'b00000000000010}; // 41, 2
    assign non_zero_info_rom[262] = {2'd2, 6'd50, 6'd51,14'b00000000100101, 14'b00000000000110}; // 37, 6
    assign non_zero_info_rom[263] = {2'd2, 6'd50, 6'd51,14'b00000000100010, 14'b00000000001001}; // 34, 9
    assign non_zero_info_rom[264] = {2'd2, 6'd50, 6'd51,14'b00000000011110, 14'b00000000001100}; // 30, 12
    assign non_zero_info_rom[265] = {2'd2, 6'd50, 6'd51,14'b00000000011011, 14'b00000000010000}; // 27, 16
    assign non_zero_info_rom[266] = {2'd2, 6'd50, 6'd51,14'b00000000010111, 14'b00000000010011}; // 23, 19
    assign non_zero_info_rom[267] = {2'd2, 6'd50, 6'd51,14'b00000000010100, 14'b00000000010110}; // 20, 22
    assign non_zero_info_rom[268] = {2'd2, 6'd50, 6'd51,14'b00000000010000, 14'b00000000011010}; // 16, 26
    assign non_zero_info_rom[269] = {2'd2, 6'd50, 6'd51,14'b00000000001101, 14'b00000000011101}; // 13, 29
    assign non_zero_info_rom[270] = {2'd2, 6'd50, 6'd51,14'b00000000001001, 14'b00000000100000}; // 9, 32
    assign non_zero_info_rom[271] = {2'd2, 6'd50, 6'd51,14'b00000000000110, 14'b00000000100100}; // 6, 36
    assign non_zero_info_rom[272] = {2'd2, 6'd50, 6'd51,14'b00000000000010, 14'b00000000100111}; // 2, 39
    assign non_zero_info_rom[273] = {2'd2, 6'd51, 6'd52,14'b00000000101000, 14'b00000000000001}; // 40, 1
    assign non_zero_info_rom[274] = {2'd2, 6'd51, 6'd52,14'b00000000100101, 14'b00000000000100}; // 37, 4
    assign non_zero_info_rom[275] = {2'd2, 6'd51, 6'd52,14'b00000000100010, 14'b00000000000111}; // 34, 7
    assign non_zero_info_rom[276] = {2'd2, 6'd51, 6'd52,14'b00000000011111, 14'b00000000001010}; // 31, 10
    assign non_zero_info_rom[277] = {2'd2, 6'd51, 6'd52,14'b00000000011100, 14'b00000000001101}; // 28, 13
    assign non_zero_info_rom[278] = {2'd2, 6'd51, 6'd52,14'b00000000011000, 14'b00000000010000}; // 24, 16
    assign non_zero_info_rom[279] = {2'd2, 6'd51, 6'd52,14'b00000000010101, 14'b00000000010011}; // 21, 19
    assign non_zero_info_rom[280] = {2'd2, 6'd51, 6'd52,14'b00000000010010, 14'b00000000010110}; // 18, 22
    assign non_zero_info_rom[281] = {2'd2, 6'd51, 6'd52,14'b00000000001111, 14'b00000000011001}; // 15, 25
    assign non_zero_info_rom[282] = {2'd2, 6'd51, 6'd52,14'b00000000001100, 14'b00000000011100}; // 12, 28
    assign non_zero_info_rom[283] = {2'd2, 6'd51, 6'd52,14'b00000000001000, 14'b00000000011111}; // 8, 31
    assign non_zero_info_rom[284] = {2'd2, 6'd51, 6'd52,14'b00000000000101, 14'b00000000100010}; // 5, 34
    assign non_zero_info_rom[285] = {2'd2, 6'd51, 6'd52,14'b00000000000010, 14'b00000000100101}; // 2, 37
    assign non_zero_info_rom[286] = {2'd2, 6'd52, 6'd53,14'b00000000100110, 14'b00000000000001}; // 38, 1
    assign non_zero_info_rom[287] = {2'd2, 6'd52, 6'd53,14'b00000000100100, 14'b00000000000100}; // 36, 4
    assign non_zero_info_rom[288] = {2'd2, 6'd52, 6'd53,14'b00000000100001, 14'b00000000000110}; // 33, 6
    assign non_zero_info_rom[289] = {2'd2, 6'd52, 6'd53,14'b00000000011110, 14'b00000000001001}; // 30, 9
    assign non_zero_info_rom[290] = {2'd2, 6'd52, 6'd53,14'b00000000011011, 14'b00000000001100}; // 27, 12
    assign non_zero_info_rom[291] = {2'd2, 6'd52, 6'd53,14'b00000000011000, 14'b00000000001111}; // 24, 15
    assign non_zero_info_rom[292] = {2'd2, 6'd52, 6'd53,14'b00000000010101, 14'b00000000010010}; // 21, 18
    assign non_zero_info_rom[293] = {2'd2, 6'd52, 6'd53,14'b00000000010010, 14'b00000000010100}; // 18, 20
    assign non_zero_info_rom[294] = {2'd2, 6'd52, 6'd53,14'b00000000001111, 14'b00000000010111}; // 15, 23
    assign non_zero_info_rom[295] = {2'd2, 6'd52, 6'd53,14'b00000000001100, 14'b00000000011010}; // 12, 26
    assign non_zero_info_rom[296] = {2'd2, 6'd52, 6'd53,14'b00000000001001, 14'b00000000011101}; // 9, 29
    assign non_zero_info_rom[297] = {2'd2, 6'd52, 6'd53,14'b00000000000111, 14'b00000000011111}; // 7, 31
    assign non_zero_info_rom[298] = {2'd2, 6'd52, 6'd53,14'b00000000000100, 14'b00000000100010}; // 4, 34
    assign non_zero_info_rom[299] = {2'd2, 6'd52, 6'd53,14'b00000000000001, 14'b00000000100101}; // 1, 37
    assign non_zero_info_rom[300] = {2'd2, 6'd53, 6'd54,14'b00000000100100, 14'b00000000000010}; // 36, 2
    assign non_zero_info_rom[301] = {2'd2, 6'd53, 6'd54,14'b00000000100001, 14'b00000000000100}; // 33, 4
    assign non_zero_info_rom[302] = {2'd2, 6'd53, 6'd54,14'b00000000011110, 14'b00000000000111}; // 30, 7
    assign non_zero_info_rom[303] = {2'd2, 6'd53, 6'd54,14'b00000000011100, 14'b00000000001001}; // 28, 9
    assign non_zero_info_rom[304] = {2'd2, 6'd53, 6'd54,14'b00000000011001, 14'b00000000001100}; // 25, 12
    assign non_zero_info_rom[305] = {2'd2, 6'd53, 6'd54,14'b00000000010110, 14'b00000000001110}; // 22, 14
    assign non_zero_info_rom[306] = {2'd2, 6'd53, 6'd54,14'b00000000010100, 14'b00000000010001}; // 20, 17
    assign non_zero_info_rom[307] = {2'd2, 6'd53, 6'd54,14'b00000000010001, 14'b00000000010100}; // 17, 20
    assign non_zero_info_rom[308] = {2'd2, 6'd53, 6'd54,14'b00000000001111, 14'b00000000010110}; // 15, 22
    assign non_zero_info_rom[309] = {2'd2, 6'd53, 6'd54,14'b00000000001100, 14'b00000000011001}; // 12, 25
    assign non_zero_info_rom[310] = {2'd2, 6'd53, 6'd54,14'b00000000001001, 14'b00000000011011}; // 9, 27
    assign non_zero_info_rom[311] = {2'd2, 6'd53, 6'd54,14'b00000000000111, 14'b00000000011110}; // 7, 30
    assign non_zero_info_rom[312] = {2'd2, 6'd53, 6'd54,14'b00000000000100, 14'b00000000100000}; // 4, 32
    assign non_zero_info_rom[313] = {2'd2, 6'd53, 6'd54,14'b00000000000001, 14'b00000000100011}; // 1, 35
    assign non_zero_info_rom[314] = {2'd2, 6'd54, 6'd55,14'b00000000100011, 14'b00000000000001}; // 35, 1
    assign non_zero_info_rom[315] = {2'd2, 6'd54, 6'd55,14'b00000000100000, 14'b00000000000011}; // 32, 3
    assign non_zero_info_rom[316] = {2'd2, 6'd54, 6'd55,14'b00000000011110, 14'b00000000000110}; // 30, 6
    assign non_zero_info_rom[317] = {2'd2, 6'd54, 6'd55,14'b00000000011100, 14'b00000000001000}; // 28, 8
    assign non_zero_info_rom[318] = {2'd2, 6'd54, 6'd55,14'b00000000011001, 14'b00000000001010}; // 25, 10
    assign non_zero_info_rom[319] = {2'd2, 6'd54, 6'd55,14'b00000000010111, 14'b00000000001101}; // 23, 13
    assign non_zero_info_rom[320] = {2'd2, 6'd54, 6'd55,14'b00000000010100, 14'b00000000001111}; // 20, 15
    assign non_zero_info_rom[321] = {2'd2, 6'd54, 6'd55,14'b00000000010010, 14'b00000000010001}; // 18, 17
    assign non_zero_info_rom[322] = {2'd2, 6'd54, 6'd55,14'b00000000010000, 14'b00000000010011}; // 16, 19
    assign non_zero_info_rom[323] = {2'd2, 6'd54, 6'd55,14'b00000000001101, 14'b00000000010110}; // 13, 22
    assign non_zero_info_rom[324] = {2'd2, 6'd54, 6'd55,14'b00000000001011, 14'b00000000011000}; // 11, 24
    assign non_zero_info_rom[325] = {2'd2, 6'd54, 6'd55,14'b00000000001000, 14'b00000000011010}; // 8, 26
    assign non_zero_info_rom[326] = {2'd2, 6'd54, 6'd55,14'b00000000000110, 14'b00000000011101}; // 6, 29
    assign non_zero_info_rom[327] = {2'd2, 6'd54, 6'd55,14'b00000000000011, 14'b00000000011111}; // 3, 31
    assign non_zero_info_rom[328] = {2'd2, 6'd54, 6'd55,14'b00000000000001, 14'b00000000100001}; // 1, 33
    assign non_zero_info_rom[329] = {2'd2, 6'd55, 6'd56,14'b00000000100001, 14'b00000000000001}; // 33, 1
    assign non_zero_info_rom[330] = {2'd2, 6'd55, 6'd56,14'b00000000011111, 14'b00000000000011}; // 31, 3
    assign non_zero_info_rom[331] = {2'd2, 6'd55, 6'd56,14'b00000000011101, 14'b00000000000101}; // 29, 5
    assign non_zero_info_rom[332] = {2'd2, 6'd55, 6'd56,14'b00000000011011, 14'b00000000000111}; // 27, 7
    assign non_zero_info_rom[333] = {2'd2, 6'd55, 6'd56,14'b00000000011000, 14'b00000000001010}; // 24, 10
    assign non_zero_info_rom[334] = {2'd2, 6'd55, 6'd56,14'b00000000010110, 14'b00000000001100}; // 22, 12
    assign non_zero_info_rom[335] = {2'd2, 6'd55, 6'd56,14'b00000000010100, 14'b00000000001110}; // 20, 14
    assign non_zero_info_rom[336] = {2'd2, 6'd55, 6'd56,14'b00000000010010, 14'b00000000010000}; // 18, 16
    assign non_zero_info_rom[337] = {2'd2, 6'd55, 6'd56,14'b00000000010000, 14'b00000000010010}; // 16, 18
    assign non_zero_info_rom[338] = {2'd2, 6'd55, 6'd56,14'b00000000001101, 14'b00000000010100}; // 13, 20
    assign non_zero_info_rom[339] = {2'd2, 6'd55, 6'd56,14'b00000000001011, 14'b00000000010110}; // 11, 22
    assign non_zero_info_rom[340] = {2'd2, 6'd55, 6'd56,14'b00000000001001, 14'b00000000011000}; // 9, 24
    assign non_zero_info_rom[341] = {2'd2, 6'd55, 6'd56,14'b00000000000111, 14'b00000000011010}; // 7, 26
    assign non_zero_info_rom[342] = {2'd2, 6'd55, 6'd56,14'b00000000000101, 14'b00000000011100}; // 5, 28
    assign non_zero_info_rom[343] = {2'd2, 6'd55, 6'd56,14'b00000000000010, 14'b00000000011110}; // 2, 30
    assign non_zero_info_rom[344] = {2'd2, 6'd55, 6'd56,14'b00000000000000, 14'b00000000100001}; // 0, 33
    assign non_zero_info_rom[345] = {2'd2, 6'd56, 6'd57,14'b00000000011111, 14'b00000000000010}; // 31, 2
    assign non_zero_info_rom[346] = {2'd2, 6'd56, 6'd57,14'b00000000011101, 14'b00000000000100}; // 29, 4
    assign non_zero_info_rom[347] = {2'd2, 6'd56, 6'd57,14'b00000000011011, 14'b00000000000110}; // 27, 6
    assign non_zero_info_rom[348] = {2'd2, 6'd56, 6'd57,14'b00000000011001, 14'b00000000000111}; // 25, 7
    assign non_zero_info_rom[349] = {2'd2, 6'd56, 6'd57,14'b00000000010111, 14'b00000000001001}; // 23, 9
    assign non_zero_info_rom[350] = {2'd2, 6'd56, 6'd57,14'b00000000010101, 14'b00000000001011}; // 21, 11
    assign non_zero_info_rom[351] = {2'd2, 6'd56, 6'd57,14'b00000000010011, 14'b00000000001101}; // 19, 13
    assign non_zero_info_rom[352] = {2'd2, 6'd56, 6'd57,14'b00000000010001, 14'b00000000001111}; // 17, 15
    assign non_zero_info_rom[353] = {2'd2, 6'd56, 6'd57,14'b00000000001111, 14'b00000000010001}; // 15, 17
    assign non_zero_info_rom[354] = {2'd2, 6'd56, 6'd57,14'b00000000001101, 14'b00000000010011}; // 13, 19
    assign non_zero_info_rom[355] = {2'd2, 6'd56, 6'd57,14'b00000000001011, 14'b00000000010101}; // 11, 21
    assign non_zero_info_rom[356] = {2'd2, 6'd56, 6'd57,14'b00000000001001, 14'b00000000010111}; // 9, 23
    assign non_zero_info_rom[357] = {2'd2, 6'd56, 6'd57,14'b00000000000111, 14'b00000000011001}; // 7, 25
    assign non_zero_info_rom[358] = {2'd2, 6'd56, 6'd57,14'b00000000000101, 14'b00000000011011}; // 5, 27
    assign non_zero_info_rom[359] = {2'd2, 6'd56, 6'd57,14'b00000000000011, 14'b00000000011100}; // 3, 28
    assign non_zero_info_rom[360] = {2'd2, 6'd56, 6'd57,14'b00000000000001, 14'b00000000011110}; // 1, 30
    assign non_zero_info_rom[361] = {2'd2, 6'd57, 6'd58,14'b00000000011110, 14'b00000000000001}; // 30, 1
    assign non_zero_info_rom[362] = {2'd2, 6'd57, 6'd58,14'b00000000011100, 14'b00000000000011}; // 28, 3
    assign non_zero_info_rom[363] = {2'd2, 6'd57, 6'd58,14'b00000000011011, 14'b00000000000100}; // 27, 4
    assign non_zero_info_rom[364] = {2'd2, 6'd57, 6'd58,14'b00000000011001, 14'b00000000000110}; // 25, 6
    assign non_zero_info_rom[365] = {2'd2, 6'd57, 6'd58,14'b00000000010111, 14'b00000000001000}; // 23, 8
    assign non_zero_info_rom[366] = {2'd2, 6'd57, 6'd58,14'b00000000010101, 14'b00000000001010}; // 21, 10
    assign non_zero_info_rom[367] = {2'd2, 6'd57, 6'd58,14'b00000000010011, 14'b00000000001011}; // 19, 11
    assign non_zero_info_rom[368] = {2'd2, 6'd57, 6'd58,14'b00000000010010, 14'b00000000001101}; // 18, 13
    assign non_zero_info_rom[369] = {2'd2, 6'd57, 6'd58,14'b00000000010000, 14'b00000000001111}; // 16, 15
    assign non_zero_info_rom[370] = {2'd2, 6'd57, 6'd58,14'b00000000001110, 14'b00000000010001}; // 14, 17
    assign non_zero_info_rom[371] = {2'd2, 6'd57, 6'd58,14'b00000000001100, 14'b00000000010010}; // 12, 18
    assign non_zero_info_rom[372] = {2'd2, 6'd57, 6'd58,14'b00000000001010, 14'b00000000010100}; // 10, 20
    assign non_zero_info_rom[373] = {2'd2, 6'd57, 6'd58,14'b00000000001000, 14'b00000000010110}; // 8, 22
    assign non_zero_info_rom[374] = {2'd2, 6'd57, 6'd58,14'b00000000000111, 14'b00000000011000}; // 7, 24
    assign non_zero_info_rom[375] = {2'd2, 6'd57, 6'd58,14'b00000000000101, 14'b00000000011001}; // 5, 25
    assign non_zero_info_rom[376] = {2'd2, 6'd57, 6'd58,14'b00000000000011, 14'b00000000011011}; // 3, 27
    assign non_zero_info_rom[377] = {2'd2, 6'd57, 6'd58,14'b00000000000001, 14'b00000000011101}; // 1, 29
    assign non_zero_info_rom[378] = {2'd2, 6'd58, 6'd59,14'b00000000011101, 14'b00000000000001}; // 29, 1
    assign non_zero_info_rom[379] = {2'd2, 6'd58, 6'd59,14'b00000000011100, 14'b00000000000010}; // 28, 2
    assign non_zero_info_rom[380] = {2'd2, 6'd58, 6'd59,14'b00000000011010, 14'b00000000000100}; // 26, 4
    assign non_zero_info_rom[381] = {2'd2, 6'd58, 6'd59,14'b00000000011000, 14'b00000000000101}; // 24, 5
    assign non_zero_info_rom[382] = {2'd2, 6'd58, 6'd59,14'b00000000010111, 14'b00000000000111}; // 23, 7
    assign non_zero_info_rom[383] = {2'd2, 6'd58, 6'd59,14'b00000000010101, 14'b00000000001001}; // 21, 9
    assign non_zero_info_rom[384] = {2'd2, 6'd58, 6'd59,14'b00000000010011, 14'b00000000001010}; // 19, 10
    assign non_zero_info_rom[385] = {2'd2, 6'd58, 6'd59,14'b00000000010010, 14'b00000000001100}; // 18, 12
    assign non_zero_info_rom[386] = {2'd2, 6'd58, 6'd59,14'b00000000010000, 14'b00000000001101}; // 16, 13
    assign non_zero_info_rom[387] = {2'd2, 6'd58, 6'd59,14'b00000000001110, 14'b00000000001111}; // 14, 15
    assign non_zero_info_rom[388] = {2'd2, 6'd58, 6'd59,14'b00000000001101, 14'b00000000010000}; // 13, 16
    assign non_zero_info_rom[389] = {2'd2, 6'd58, 6'd59,14'b00000000001011, 14'b00000000010010}; // 11, 18
    assign non_zero_info_rom[390] = {2'd2, 6'd58, 6'd59,14'b00000000001001, 14'b00000000010100}; // 9, 20
    assign non_zero_info_rom[391] = {2'd2, 6'd58, 6'd59,14'b00000000001000, 14'b00000000010101}; // 8, 21
    assign non_zero_info_rom[392] = {2'd2, 6'd58, 6'd59,14'b00000000000110, 14'b00000000010111}; // 6, 23
    assign non_zero_info_rom[393] = {2'd2, 6'd58, 6'd59,14'b00000000000100, 14'b00000000011000}; // 4, 24
    assign non_zero_info_rom[394] = {2'd2, 6'd58, 6'd59,14'b00000000000011, 14'b00000000011010}; // 3, 26
    assign non_zero_info_rom[395] = {2'd2, 6'd58, 6'd59,14'b00000000000001, 14'b00000000011100}; // 1, 28
    assign non_zero_info_rom[396] = {2'd2, 6'd59, 6'd60,14'b00000000011100, 14'b00000000000001}; // 28, 1
    assign non_zero_info_rom[397] = {2'd2, 6'd59, 6'd60,14'b00000000011010, 14'b00000000000010}; // 26, 2
    assign non_zero_info_rom[398] = {2'd2, 6'd59, 6'd60,14'b00000000011001, 14'b00000000000011}; // 25, 3
    assign non_zero_info_rom[399] = {2'd2, 6'd59, 6'd60,14'b00000000010111, 14'b00000000000101}; // 23, 5
    assign non_zero_info_rom[400] = {2'd2, 6'd59, 6'd60,14'b00000000010110, 14'b00000000000110}; // 22, 6
    assign non_zero_info_rom[401] = {2'd2, 6'd59, 6'd60,14'b00000000010100, 14'b00000000001000}; // 20, 8
    assign non_zero_info_rom[402] = {2'd2, 6'd59, 6'd60,14'b00000000010011, 14'b00000000001001}; // 19, 9
    assign non_zero_info_rom[403] = {2'd2, 6'd59, 6'd60,14'b00000000010001, 14'b00000000001011}; // 17, 11
    assign non_zero_info_rom[404] = {2'd2, 6'd59, 6'd60,14'b00000000010000, 14'b00000000001100}; // 16, 12
    assign non_zero_info_rom[405] = {2'd2, 6'd59, 6'd60,14'b00000000001110, 14'b00000000001110}; // 14, 14
    assign non_zero_info_rom[406] = {2'd2, 6'd59, 6'd60,14'b00000000001101, 14'b00000000001111}; // 13, 15
    assign non_zero_info_rom[407] = {2'd2, 6'd59, 6'd60,14'b00000000001011, 14'b00000000010000}; // 11, 16
    assign non_zero_info_rom[408] = {2'd2, 6'd59, 6'd60,14'b00000000001010, 14'b00000000010010}; // 10, 18
    assign non_zero_info_rom[409] = {2'd2, 6'd59, 6'd60,14'b00000000001000, 14'b00000000010011}; // 8, 19
    assign non_zero_info_rom[410] = {2'd2, 6'd59, 6'd60,14'b00000000000111, 14'b00000000010101}; // 7, 21
    assign non_zero_info_rom[411] = {2'd2, 6'd59, 6'd60,14'b00000000000101, 14'b00000000010110}; // 5, 22
    assign non_zero_info_rom[412] = {2'd2, 6'd59, 6'd60,14'b00000000000100, 14'b00000000011000}; // 4, 24
    assign non_zero_info_rom[413] = {2'd2, 6'd59, 6'd60,14'b00000000000010, 14'b00000000011001}; // 2, 25
    assign non_zero_info_rom[414] = {2'd2, 6'd59, 6'd60,14'b00000000000001, 14'b00000000011011}; // 1, 27
    assign non_zero_info_rom[415] = {2'd2, 6'd60, 6'd61,14'b00000000011010, 14'b00000000000001}; // 26, 1
    assign non_zero_info_rom[416] = {2'd2, 6'd60, 6'd61,14'b00000000011001, 14'b00000000000010}; // 25, 2
    assign non_zero_info_rom[417] = {2'd2, 6'd60, 6'd61,14'b00000000011000, 14'b00000000000011}; // 24, 3
    assign non_zero_info_rom[418] = {2'd2, 6'd60, 6'd61,14'b00000000010110, 14'b00000000000101}; // 22, 5
    assign non_zero_info_rom[419] = {2'd2, 6'd60, 6'd61,14'b00000000010101, 14'b00000000000110}; // 21, 6
    assign non_zero_info_rom[420] = {2'd2, 6'd60, 6'd61,14'b00000000010100, 14'b00000000000111}; // 20, 7
    assign non_zero_info_rom[421] = {2'd2, 6'd60, 6'd61,14'b00000000010010, 14'b00000000001001}; // 18, 9
    assign non_zero_info_rom[422] = {2'd2, 6'd60, 6'd61,14'b00000000010001, 14'b00000000001010}; // 17, 10
    assign non_zero_info_rom[423] = {2'd2, 6'd60, 6'd61,14'b00000000001111, 14'b00000000001011}; // 15, 11
    assign non_zero_info_rom[424] = {2'd2, 6'd60, 6'd61,14'b00000000001110, 14'b00000000001101}; // 14, 13
    assign non_zero_info_rom[425] = {2'd2, 6'd60, 6'd61,14'b00000000001101, 14'b00000000001110}; // 13, 14
    assign non_zero_info_rom[426] = {2'd2, 6'd60, 6'd61,14'b00000000001011, 14'b00000000001111}; // 11, 15
    assign non_zero_info_rom[427] = {2'd2, 6'd60, 6'd61,14'b00000000001010, 14'b00000000010001}; // 10, 17
    assign non_zero_info_rom[428] = {2'd2, 6'd60, 6'd61,14'b00000000001001, 14'b00000000010010}; // 9, 18
    assign non_zero_info_rom[429] = {2'd2, 6'd60, 6'd61,14'b00000000000111, 14'b00000000010011}; // 7, 19
    assign non_zero_info_rom[430] = {2'd2, 6'd60, 6'd61,14'b00000000000110, 14'b00000000010100}; // 6, 20
    assign non_zero_info_rom[431] = {2'd2, 6'd60, 6'd61,14'b00000000000100, 14'b00000000010110}; // 4, 22
    assign non_zero_info_rom[432] = {2'd2, 6'd60, 6'd61,14'b00000000000011, 14'b00000000010111}; // 3, 23
    assign non_zero_info_rom[433] = {2'd2, 6'd60, 6'd61,14'b00000000000010, 14'b00000000011000}; // 2, 24
    assign non_zero_info_rom[434] = {2'd2, 6'd60, 6'd61,14'b00000000000000, 14'b00000000011010}; // 0, 26
    assign non_zero_info_rom[435] = {2'd2, 6'd61, 6'd62,14'b00000000011001, 14'b00000000000001}; // 25, 1
    assign non_zero_info_rom[436] = {2'd2, 6'd61, 6'd62,14'b00000000011000, 14'b00000000000010}; // 24, 2
    assign non_zero_info_rom[437] = {2'd2, 6'd61, 6'd62,14'b00000000010110, 14'b00000000000011}; // 22, 3
    assign non_zero_info_rom[438] = {2'd2, 6'd61, 6'd62,14'b00000000010101, 14'b00000000000101}; // 21, 5
    assign non_zero_info_rom[439] = {2'd2, 6'd61, 6'd62,14'b00000000010100, 14'b00000000000110}; // 20, 6
    assign non_zero_info_rom[440] = {2'd2, 6'd61, 6'd62,14'b00000000010011, 14'b00000000000111}; // 19, 7
    assign non_zero_info_rom[441] = {2'd2, 6'd61, 6'd62,14'b00000000010001, 14'b00000000001000}; // 17, 8
    assign non_zero_info_rom[442] = {2'd2, 6'd61, 6'd62,14'b00000000010000, 14'b00000000001001}; // 16, 9
    assign non_zero_info_rom[443] = {2'd2, 6'd61, 6'd62,14'b00000000001111, 14'b00000000001011}; // 15, 11
    assign non_zero_info_rom[444] = {2'd2, 6'd61, 6'd62,14'b00000000001110, 14'b00000000001100}; // 14, 12
    assign non_zero_info_rom[445] = {2'd2, 6'd61, 6'd62,14'b00000000001100, 14'b00000000001101}; // 12, 13
    assign non_zero_info_rom[446] = {2'd2, 6'd61, 6'd62,14'b00000000001011, 14'b00000000001110}; // 11, 14
    assign non_zero_info_rom[447] = {2'd2, 6'd61, 6'd62,14'b00000000001010, 14'b00000000001111}; // 10, 15
    assign non_zero_info_rom[448] = {2'd2, 6'd61, 6'd62,14'b00000000001001, 14'b00000000010001}; // 9, 17
    assign non_zero_info_rom[449] = {2'd2, 6'd61, 6'd62,14'b00000000000111, 14'b00000000010010}; // 7, 18
    assign non_zero_info_rom[450] = {2'd2, 6'd61, 6'd62,14'b00000000000110, 14'b00000000010011}; // 6, 19
    assign non_zero_info_rom[451] = {2'd2, 6'd61, 6'd62,14'b00000000000101, 14'b00000000010100}; // 5, 20
    assign non_zero_info_rom[452] = {2'd2, 6'd61, 6'd62,14'b00000000000100, 14'b00000000010101}; // 4, 21
    assign non_zero_info_rom[453] = {2'd2, 6'd61, 6'd62,14'b00000000000010, 14'b00000000010111}; // 2, 23
    assign non_zero_info_rom[454] = {2'd2, 6'd61, 6'd62,14'b00000000000001, 14'b00000000011000}; // 1, 24
    assign non_zero_info_rom[455] = {2'd2, 6'd62, 6'd63,14'b00000000011001, 14'b00000000000000}; // 25, 0
    assign non_zero_info_rom[456] = {2'd2, 6'd62, 6'd63,14'b00000000010111, 14'b00000000000001}; // 23, 1
    assign non_zero_info_rom[457] = {2'd2, 6'd62, 6'd63,14'b00000000010110, 14'b00000000000010}; // 22, 2
    assign non_zero_info_rom[458] = {2'd2, 6'd62, 6'd63,14'b00000000010101, 14'b00000000000011}; // 21, 3
    assign non_zero_info_rom[459] = {2'd2, 6'd62, 6'd63,14'b00000000010100, 14'b00000000000101}; // 20, 5
    assign non_zero_info_rom[460] = {2'd2, 6'd62, 6'd63,14'b00000000010011, 14'b00000000000110}; // 19, 6
    assign non_zero_info_rom[461] = {2'd2, 6'd62, 6'd63,14'b00000000010010, 14'b00000000000111}; // 18, 7
    assign non_zero_info_rom[462] = {2'd2, 6'd62, 6'd63,14'b00000000010001, 14'b00000000001000}; // 17, 8
    assign non_zero_info_rom[463] = {2'd2, 6'd62, 6'd63,14'b00000000001111, 14'b00000000001001}; // 15, 9
    assign non_zero_info_rom[464] = {2'd2, 6'd62, 6'd63,14'b00000000001110, 14'b00000000001010}; // 14, 10
    assign non_zero_info_rom[465] = {2'd2, 6'd62, 6'd63,14'b00000000001101, 14'b00000000001011}; // 13, 11
    assign non_zero_info_rom[466] = {2'd2, 6'd62, 6'd63,14'b00000000001100, 14'b00000000001100}; // 12, 12
    assign non_zero_info_rom[467] = {2'd2, 6'd62, 6'd63,14'b00000000001011, 14'b00000000001101}; // 11, 13
    assign non_zero_info_rom[468] = {2'd2, 6'd62, 6'd63,14'b00000000001010, 14'b00000000001110}; // 10, 14
    assign non_zero_info_rom[469] = {2'd2, 6'd62, 6'd63,14'b00000000001001, 14'b00000000001111}; // 9, 15
    assign non_zero_info_rom[470] = {2'd2, 6'd62, 6'd63,14'b00000000000111, 14'b00000000010001}; // 7, 17
    assign non_zero_info_rom[471] = {2'd2, 6'd62, 6'd63,14'b00000000000110, 14'b00000000010010}; // 6, 18
    assign non_zero_info_rom[472] = {2'd2, 6'd62, 6'd63,14'b00000000000101, 14'b00000000010011}; // 5, 19
    assign non_zero_info_rom[473] = {2'd2, 6'd62, 6'd63,14'b00000000000100, 14'b00000000010100}; // 4, 20
    assign non_zero_info_rom[474] = {2'd2, 6'd62, 6'd63,14'b00000000000011, 14'b00000000010101}; // 3, 21
    assign non_zero_info_rom[475] = {2'd2, 6'd62, 6'd63,14'b00000000000010, 14'b00000000010110}; // 2, 22
    assign non_zero_info_rom[476] = {2'd2, 6'd62, 6'd63,14'b00000000000001, 14'b00000000010111}; // 1, 23
    assign non_zero_info_rom[477] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010111, 14'bxxxxxxxxxxxxxx}; // 23
    assign non_zero_info_rom[478] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010110, 14'bxxxxxxxxxxxxxx}; // 22
    assign non_zero_info_rom[479] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010101, 14'bxxxxxxxxxxxxxx}; // 21
    assign non_zero_info_rom[480] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010100, 14'bxxxxxxxxxxxxxx}; // 20
    assign non_zero_info_rom[481] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010011, 14'bxxxxxxxxxxxxxx}; // 19
    assign non_zero_info_rom[482] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010010, 14'bxxxxxxxxxxxxxx}; // 18
    assign non_zero_info_rom[483] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010001, 14'bxxxxxxxxxxxxxx}; // 17
    assign non_zero_info_rom[484] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000010000, 14'bxxxxxxxxxxxxxx}; // 16
    assign non_zero_info_rom[485] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001111, 14'bxxxxxxxxxxxxxx}; // 15
    assign non_zero_info_rom[486] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001110, 14'bxxxxxxxxxxxxxx}; // 14
    assign non_zero_info_rom[487] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001101, 14'bxxxxxxxxxxxxxx}; // 13
    assign non_zero_info_rom[488] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001100, 14'bxxxxxxxxxxxxxx}; // 12
    assign non_zero_info_rom[489] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001011, 14'bxxxxxxxxxxxxxx}; // 11
    assign non_zero_info_rom[490] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001010, 14'bxxxxxxxxxxxxxx}; // 10
    assign non_zero_info_rom[491] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001001, 14'bxxxxxxxxxxxxxx}; // 9
    assign non_zero_info_rom[492] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000001000, 14'bxxxxxxxxxxxxxx}; // 8
    assign non_zero_info_rom[493] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000110, 14'bxxxxxxxxxxxxxx}; // 6
    assign non_zero_info_rom[494] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000101, 14'bxxxxxxxxxxxxxx}; // 5
    assign non_zero_info_rom[495] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000100, 14'bxxxxxxxxxxxxxx}; // 4
    assign non_zero_info_rom[496] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000011, 14'bxxxxxxxxxxxxxx}; // 3
    assign non_zero_info_rom[497] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000010, 14'bxxxxxxxxxxxxxx}; // 2
    assign non_zero_info_rom[498] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000001, 14'bxxxxxxxxxxxxxx}; // 1
    assign non_zero_info_rom[499] = {2'd1, 6'd63, 6'bxxxxxx,14'b00000000000000, 14'bxxxxxxxxxxxxxx}; // 0
    assign non_zero_info_rom[500] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[501] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[502] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[503] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[504] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[505] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[506] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[507] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[508] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[509] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[510] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[511] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 
    assign non_zero_info_rom[512] = {2'd0, 6'bxxxxxx, 6'bxxxxxx,14'bxxxxxxxxxxxxxx, 14'bxxxxxxxxxxxxxx}; // 

endmodule