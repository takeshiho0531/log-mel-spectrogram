module hann_window_rom (
    input clk,
    input rst,
    input [9:0] window_num,
    output [13:0] window_coef
  );
    wire signed [13:0] window_rom[0:1023];
    
    assign window_coef = window_rom[window_num];

    assign window_rom[0]={1'b0, 13'd0};
    assign window_rom[1]={1'b0, 13'd0};
    assign window_rom[2]={1'b0, 13'd0};
    assign window_rom[3]={1'b0, 13'd1};
    assign window_rom[4]={1'b0, 13'd1};
    assign window_rom[5]={1'b0, 13'd2};
    assign window_rom[6]={1'b0, 13'd3};
    assign window_rom[7]={1'b0, 13'd4};
    assign window_rom[8]={1'b0, 13'd5};
    assign window_rom[9]={1'b0, 13'd6};
    assign window_rom[10]={1'b0, 13'd8};
    assign window_rom[11]={1'b0, 13'd9};
    assign window_rom[12]={1'b0, 13'd11};
    assign window_rom[13]={1'b0, 13'd13};
    assign window_rom[14]={1'b0, 13'd15};
    assign window_rom[15]={1'b0, 13'd17};
    assign window_rom[16]={1'b0, 13'd20};
    assign window_rom[17]={1'b0, 13'd22};
    assign window_rom[18]={1'b0, 13'd25};
    assign window_rom[19]={1'b0, 13'd28};
    assign window_rom[20]={1'b0, 13'd30};
    assign window_rom[21]={1'b0, 13'd34};
    assign window_rom[22]={1'b0, 13'd37};
    assign window_rom[23]={1'b0, 13'd40};
    assign window_rom[24]={1'b0, 13'd44};
    assign window_rom[25]={1'b0, 13'd48};
    assign window_rom[26]={1'b0, 13'd51};
    assign window_rom[27]={1'b0, 13'd56};
    assign window_rom[28]={1'b0, 13'd60};
    assign window_rom[29]={1'b0, 13'd64};
    assign window_rom[30]={1'b0, 13'd69};
    assign window_rom[31]={1'b0, 13'd73};
    assign window_rom[32]={1'b0, 13'd78};
    assign window_rom[33]={1'b0, 13'd83};
    assign window_rom[34]={1'b0, 13'd88};
    assign window_rom[35]={1'b0, 13'd93};
    assign window_rom[36]={1'b0, 13'd99};
    assign window_rom[37]={1'b0, 13'd104};
    assign window_rom[38]={1'b0, 13'd110};
    assign window_rom[39]={1'b0, 13'd116};
    assign window_rom[40]={1'b0, 13'd122};
    assign window_rom[41]={1'b0, 13'd128};
    assign window_rom[42]={1'b0, 13'd134};
    assign window_rom[43]={1'b0, 13'd140};
    assign window_rom[44]={1'b0, 13'd147};
    assign window_rom[45]={1'b0, 13'd154};
    assign window_rom[46]={1'b0, 13'd160};
    assign window_rom[47]={1'b0, 13'd167};
    assign window_rom[48]={1'b0, 13'd175};
    assign window_rom[49]={1'b0, 13'd182};
    assign window_rom[50]={1'b0, 13'd189};
    assign window_rom[51]={1'b0, 13'd197};
    assign window_rom[52]={1'b0, 13'd205};
    assign window_rom[53]={1'b0, 13'd213};
    assign window_rom[54]={1'b0, 13'd221};
    assign window_rom[55]={1'b0, 13'd229};
    assign window_rom[56]={1'b0, 13'd237};
    assign window_rom[57]={1'b0, 13'd245};
    assign window_rom[58]={1'b0, 13'd254};
    assign window_rom[59]={1'b0, 13'd263};
    assign window_rom[60]={1'b0, 13'd272};
    assign window_rom[61]={1'b0, 13'd281};
    assign window_rom[62]={1'b0, 13'd290};
    assign window_rom[63]={1'b0, 13'd299};
    assign window_rom[64]={1'b0, 13'd309};
    assign window_rom[65]={1'b0, 13'd318};
    assign window_rom[66]={1'b0, 13'd328};
    assign window_rom[67]={1'b0, 13'd338};
    assign window_rom[68]={1'b0, 13'd348};
    assign window_rom[69]={1'b0, 13'd358};
    assign window_rom[70]={1'b0, 13'd368};
    assign window_rom[71]={1'b0, 13'd379};
    assign window_rom[72]={1'b0, 13'd389};
    assign window_rom[73]={1'b0, 13'd400};
    assign window_rom[74]={1'b0, 13'd411};
    assign window_rom[75]={1'b0, 13'd422};
    assign window_rom[76]={1'b0, 13'd433};
    assign window_rom[77]={1'b0, 13'd444};
    assign window_rom[78]={1'b0, 13'd456};
    assign window_rom[79]={1'b0, 13'd467};
    assign window_rom[80]={1'b0, 13'd479};
    assign window_rom[81]={1'b0, 13'd491};
    assign window_rom[82]={1'b0, 13'd503};
    assign window_rom[83]={1'b0, 13'd515};
    assign window_rom[84]={1'b0, 13'd527};
    assign window_rom[85]={1'b0, 13'd539};
    assign window_rom[86]={1'b0, 13'd552};
    assign window_rom[87]={1'b0, 13'd564};
    assign window_rom[88]={1'b0, 13'd577};
    assign window_rom[89]={1'b0, 13'd590};
    assign window_rom[90]={1'b0, 13'd603};
    assign window_rom[91]={1'b0, 13'd616};
    assign window_rom[92]={1'b0, 13'd629};
    assign window_rom[93]={1'b0, 13'd643};
    assign window_rom[94]={1'b0, 13'd656};
    assign window_rom[95]={1'b0, 13'd670};
    assign window_rom[96]={1'b0, 13'd683};
    assign window_rom[97]={1'b0, 13'd697};
    assign window_rom[98]={1'b0, 13'd711};
    assign window_rom[99]={1'b0, 13'd725};
    assign window_rom[100]={1'b0, 13'd740};
    assign window_rom[101]={1'b0, 13'd754};
    assign window_rom[102]={1'b0, 13'd769};
    assign window_rom[103]={1'b0, 13'd783};
    assign window_rom[104]={1'b0, 13'd798};
    assign window_rom[105]={1'b0, 13'd813};
    assign window_rom[106]={1'b0, 13'd828};
    assign window_rom[107]={1'b0, 13'd843};
    assign window_rom[108]={1'b0, 13'd858};
    assign window_rom[109]={1'b0, 13'd874};
    assign window_rom[110]={1'b0, 13'd889};
    assign window_rom[111]={1'b0, 13'd905};
    assign window_rom[112]={1'b0, 13'd920};
    assign window_rom[113]={1'b0, 13'd936};
    assign window_rom[114]={1'b0, 13'd952};
    assign window_rom[115]={1'b0, 13'd968};
    assign window_rom[116]={1'b0, 13'd985};
    assign window_rom[117]={1'b0, 13'd1001};
    assign window_rom[118]={1'b0, 13'd1017};
    assign window_rom[119]={1'b0, 13'd1034};
    assign window_rom[120]={1'b0, 13'd1050};
    assign window_rom[121]={1'b0, 13'd1067};
    assign window_rom[122]={1'b0, 13'd1084};
    assign window_rom[123]={1'b0, 13'd1101};
    assign window_rom[124]={1'b0, 13'd1118};
    assign window_rom[125]={1'b0, 13'd1135};
    assign window_rom[126]={1'b0, 13'd1153};
    assign window_rom[127]={1'b0, 13'd1170};
    assign window_rom[128]={1'b0, 13'd1188};
    assign window_rom[129]={1'b0, 13'd1205};
    assign window_rom[130]={1'b0, 13'd1223};
    assign window_rom[131]={1'b0, 13'd1241};
    assign window_rom[132]={1'b0, 13'd1259};
    assign window_rom[133]={1'b0, 13'd1277};
    assign window_rom[134]={1'b0, 13'd1295};
    assign window_rom[135]={1'b0, 13'd1313};
    assign window_rom[136]={1'b0, 13'd1332};
    assign window_rom[137]={1'b0, 13'd1350};
    assign window_rom[138]={1'b0, 13'd1369};
    assign window_rom[139]={1'b0, 13'd1388};
    assign window_rom[140]={1'b0, 13'd1406};
    assign window_rom[141]={1'b0, 13'd1425};
    assign window_rom[142]={1'b0, 13'd1444};
    assign window_rom[143]={1'b0, 13'd1463};
    assign window_rom[144]={1'b0, 13'd1483};
    assign window_rom[145]={1'b0, 13'd1502};
    assign window_rom[146]={1'b0, 13'd1521};
    assign window_rom[147]={1'b0, 13'd1541};
    assign window_rom[148]={1'b0, 13'd1560};
    assign window_rom[149]={1'b0, 13'd1580};
    assign window_rom[150]={1'b0, 13'd1600};
    assign window_rom[151]={1'b0, 13'd1620};
    assign window_rom[152]={1'b0, 13'd1639};
    assign window_rom[153]={1'b0, 13'd1659};
    assign window_rom[154]={1'b0, 13'd1680};
    assign window_rom[155]={1'b0, 13'd1700};
    assign window_rom[156]={1'b0, 13'd1720};
    assign window_rom[157]={1'b0, 13'd1741};
    assign window_rom[158]={1'b0, 13'd1761};
    assign window_rom[159]={1'b0, 13'd1782};
    assign window_rom[160]={1'b0, 13'd1802};
    assign window_rom[161]={1'b0, 13'd1823};
    assign window_rom[162]={1'b0, 13'd1844};
    assign window_rom[163]={1'b0, 13'd1865};
    assign window_rom[164]={1'b0, 13'd1886};
    assign window_rom[165]={1'b0, 13'd1907};
    assign window_rom[166]={1'b0, 13'd1928};
    assign window_rom[167]={1'b0, 13'd1949};
    assign window_rom[168]={1'b0, 13'd1970};
    assign window_rom[169]={1'b0, 13'd1992};
    assign window_rom[170]={1'b0, 13'd2013};
    assign window_rom[171]={1'b0, 13'd2035};
    assign window_rom[172]={1'b0, 13'd2056};
    assign window_rom[173]={1'b0, 13'd2078};
    assign window_rom[174]={1'b0, 13'd2100};
    assign window_rom[175]={1'b0, 13'd2122};
    assign window_rom[176]={1'b0, 13'd2144};
    assign window_rom[177]={1'b0, 13'd2165};
    assign window_rom[178]={1'b0, 13'd2188};
    assign window_rom[179]={1'b0, 13'd2210};
    assign window_rom[180]={1'b0, 13'd2232};
    assign window_rom[181]={1'b0, 13'd2254};
    assign window_rom[182]={1'b0, 13'd2276};
    assign window_rom[183]={1'b0, 13'd2299};
    assign window_rom[184]={1'b0, 13'd2321};
    assign window_rom[185]={1'b0, 13'd2344};
    assign window_rom[186]={1'b0, 13'd2366};
    assign window_rom[187]={1'b0, 13'd2389};
    assign window_rom[188]={1'b0, 13'd2412};
    assign window_rom[189]={1'b0, 13'd2435};
    assign window_rom[190]={1'b0, 13'd2457};
    assign window_rom[191]={1'b0, 13'd2480};
    assign window_rom[192]={1'b0, 13'd2503};
    assign window_rom[193]={1'b0, 13'd2526};
    assign window_rom[194]={1'b0, 13'd2549};
    assign window_rom[195]={1'b0, 13'd2572};
    assign window_rom[196]={1'b0, 13'd2596};
    assign window_rom[197]={1'b0, 13'd2619};
    assign window_rom[198]={1'b0, 13'd2642};
    assign window_rom[199]={1'b0, 13'd2666};
    assign window_rom[200]={1'b0, 13'd2689};
    assign window_rom[201]={1'b0, 13'd2712};
    assign window_rom[202]={1'b0, 13'd2736};
    assign window_rom[203]={1'b0, 13'd2759};
    assign window_rom[204]={1'b0, 13'd2783};
    assign window_rom[205]={1'b0, 13'd2807};
    assign window_rom[206]={1'b0, 13'd2830};
    assign window_rom[207]={1'b0, 13'd2854};
    assign window_rom[208]={1'b0, 13'd2878};
    assign window_rom[209]={1'b0, 13'd2902};
    assign window_rom[210]={1'b0, 13'd2926};
    assign window_rom[211]={1'b0, 13'd2950};
    assign window_rom[212]={1'b0, 13'd2974};
    assign window_rom[213]={1'b0, 13'd2998};
    assign window_rom[214]={1'b0, 13'd3022};
    assign window_rom[215]={1'b0, 13'd3046};
    assign window_rom[216]={1'b0, 13'd3070};
    assign window_rom[217]={1'b0, 13'd3094};
    assign window_rom[218]={1'b0, 13'd3118};
    assign window_rom[219]={1'b0, 13'd3142};
    assign window_rom[220]={1'b0, 13'd3167};
    assign window_rom[221]={1'b0, 13'd3191};
    assign window_rom[222]={1'b0, 13'd3215};
    assign window_rom[223]={1'b0, 13'd3240};
    assign window_rom[224]={1'b0, 13'd3264};
    assign window_rom[225]={1'b0, 13'd3288};
    assign window_rom[226]={1'b0, 13'd3313};
    assign window_rom[227]={1'b0, 13'd3337};
    assign window_rom[228]={1'b0, 13'd3362};
    assign window_rom[229]={1'b0, 13'd3386};
    assign window_rom[230]={1'b0, 13'd3411};
    assign window_rom[231]={1'b0, 13'd3435};
    assign window_rom[232]={1'b0, 13'd3460};
    assign window_rom[233]={1'b0, 13'd3485};
    assign window_rom[234]={1'b0, 13'd3509};
    assign window_rom[235]={1'b0, 13'd3534};
    assign window_rom[236]={1'b0, 13'd3559};
    assign window_rom[237]={1'b0, 13'd3583};
    assign window_rom[238]={1'b0, 13'd3608};
    assign window_rom[239]={1'b0, 13'd3633};
    assign window_rom[240]={1'b0, 13'd3658};
    assign window_rom[241]={1'b0, 13'd3682};
    assign window_rom[242]={1'b0, 13'd3707};
    assign window_rom[243]={1'b0, 13'd3732};
    assign window_rom[244]={1'b0, 13'd3757};
    assign window_rom[245]={1'b0, 13'd3782};
    assign window_rom[246]={1'b0, 13'd3806};
    assign window_rom[247]={1'b0, 13'd3831};
    assign window_rom[248]={1'b0, 13'd3856};
    assign window_rom[249]={1'b0, 13'd3881};
    assign window_rom[250]={1'b0, 13'd3906};
    assign window_rom[251]={1'b0, 13'd3931};
    assign window_rom[252]={1'b0, 13'd3956};
    assign window_rom[253]={1'b0, 13'd3980};
    assign window_rom[254]={1'b0, 13'd4005};
    assign window_rom[255]={1'b0, 13'd4030};
    assign window_rom[256]={1'b0, 13'd4055};
    assign window_rom[257]={1'b0, 13'd4080};
    assign window_rom[258]={1'b0, 13'd4105};
    assign window_rom[259]={1'b0, 13'd4130};
    assign window_rom[260]={1'b0, 13'd4155};
    assign window_rom[261]={1'b0, 13'd4179};
    assign window_rom[262]={1'b0, 13'd4204};
    assign window_rom[263]={1'b0, 13'd4229};
    assign window_rom[264]={1'b0, 13'd4254};
    assign window_rom[265]={1'b0, 13'd4279};
    assign window_rom[266]={1'b0, 13'd4304};
    assign window_rom[267]={1'b0, 13'd4329};
    assign window_rom[268]={1'b0, 13'd4353};
    assign window_rom[269]={1'b0, 13'd4378};
    assign window_rom[270]={1'b0, 13'd4403};
    assign window_rom[271]={1'b0, 13'd4428};
    assign window_rom[272]={1'b0, 13'd4453};
    assign window_rom[273]={1'b0, 13'd4477};
    assign window_rom[274]={1'b0, 13'd4502};
    assign window_rom[275]={1'b0, 13'd4527};
    assign window_rom[276]={1'b0, 13'd4551};
    assign window_rom[277]={1'b0, 13'd4576};
    assign window_rom[278]={1'b0, 13'd4601};
    assign window_rom[279]={1'b0, 13'd4625};
    assign window_rom[280]={1'b0, 13'd4650};
    assign window_rom[281]={1'b0, 13'd4675};
    assign window_rom[282]={1'b0, 13'd4699};
    assign window_rom[283]={1'b0, 13'd4724};
    assign window_rom[284]={1'b0, 13'd4748};
    assign window_rom[285]={1'b0, 13'd4773};
    assign window_rom[286]={1'b0, 13'd4797};
    assign window_rom[287]={1'b0, 13'd4822};
    assign window_rom[288]={1'b0, 13'd4846};
    assign window_rom[289]={1'b0, 13'd4871};
    assign window_rom[290]={1'b0, 13'd4895};
    assign window_rom[291]={1'b0, 13'd4919};
    assign window_rom[292]={1'b0, 13'd4944};
    assign window_rom[293]={1'b0, 13'd4968};
    assign window_rom[294]={1'b0, 13'd4992};
    assign window_rom[295]={1'b0, 13'd5016};
    assign window_rom[296]={1'b0, 13'd5040};
    assign window_rom[297]={1'b0, 13'd5064};
    assign window_rom[298]={1'b0, 13'd5089};
    assign window_rom[299]={1'b0, 13'd5113};
    assign window_rom[300]={1'b0, 13'd5137};
    assign window_rom[301]={1'b0, 13'd5161};
    assign window_rom[302]={1'b0, 13'd5184};
    assign window_rom[303]={1'b0, 13'd5208};
    assign window_rom[304]={1'b0, 13'd5232};
    assign window_rom[305]={1'b0, 13'd5256};
    assign window_rom[306]={1'b0, 13'd5280};
    assign window_rom[307]={1'b0, 13'd5303};
    assign window_rom[308]={1'b0, 13'd5327};
    assign window_rom[309]={1'b0, 13'd5351};
    assign window_rom[310]={1'b0, 13'd5374};
    assign window_rom[311]={1'b0, 13'd5398};
    assign window_rom[312]={1'b0, 13'd5421};
    assign window_rom[313]={1'b0, 13'd5445};
    assign window_rom[314]={1'b0, 13'd5468};
    assign window_rom[315]={1'b0, 13'd5491};
    assign window_rom[316]={1'b0, 13'd5514};
    assign window_rom[317]={1'b0, 13'd5538};
    assign window_rom[318]={1'b0, 13'd5561};
    assign window_rom[319]={1'b0, 13'd5584};
    assign window_rom[320]={1'b0, 13'd5607};
    assign window_rom[321]={1'b0, 13'd5630};
    assign window_rom[322]={1'b0, 13'd5653};
    assign window_rom[323]={1'b0, 13'd5676};
    assign window_rom[324]={1'b0, 13'd5698};
    assign window_rom[325]={1'b0, 13'd5721};
    assign window_rom[326]={1'b0, 13'd5744};
    assign window_rom[327]={1'b0, 13'd5766};
    assign window_rom[328]={1'b0, 13'd5789};
    assign window_rom[329]={1'b0, 13'd5811};
    assign window_rom[330]={1'b0, 13'd5834};
    assign window_rom[331]={1'b0, 13'd5856};
    assign window_rom[332]={1'b0, 13'd5878};
    assign window_rom[333]={1'b0, 13'd5900};
    assign window_rom[334]={1'b0, 13'd5923};
    assign window_rom[335]={1'b0, 13'd5945};
    assign window_rom[336]={1'b0, 13'd5967};
    assign window_rom[337]={1'b0, 13'd5988};
    assign window_rom[338]={1'b0, 13'd6010};
    assign window_rom[339]={1'b0, 13'd6032};
    assign window_rom[340]={1'b0, 13'd6054};
    assign window_rom[341]={1'b0, 13'd6075};
    assign window_rom[342]={1'b0, 13'd6097};
    assign window_rom[343]={1'b0, 13'd6118};
    assign window_rom[344]={1'b0, 13'd6140};
    assign window_rom[345]={1'b0, 13'd6161};
    assign window_rom[346]={1'b0, 13'd6182};
    assign window_rom[347]={1'b0, 13'd6203};
    assign window_rom[348]={1'b0, 13'd6224};
    assign window_rom[349]={1'b0, 13'd6245};
    assign window_rom[350]={1'b0, 13'd6266};
    assign window_rom[351]={1'b0, 13'd6287};
    assign window_rom[352]={1'b0, 13'd6308};
    assign window_rom[353]={1'b0, 13'd6329};
    assign window_rom[354]={1'b0, 13'd6349};
    assign window_rom[355]={1'b0, 13'd6370};
    assign window_rom[356]={1'b0, 13'd6390};
    assign window_rom[357]={1'b0, 13'd6410};
    assign window_rom[358]={1'b0, 13'd6430};
    assign window_rom[359]={1'b0, 13'd6451};
    assign window_rom[360]={1'b0, 13'd6471};
    assign window_rom[361]={1'b0, 13'd6491};
    assign window_rom[362]={1'b0, 13'd6510};
    assign window_rom[363]={1'b0, 13'd6530};
    assign window_rom[364]={1'b0, 13'd6550};
    assign window_rom[365]={1'b0, 13'd6569};
    assign window_rom[366]={1'b0, 13'd6589};
    assign window_rom[367]={1'b0, 13'd6608};
    assign window_rom[368]={1'b0, 13'd6628};
    assign window_rom[369]={1'b0, 13'd6647};
    assign window_rom[370]={1'b0, 13'd6666};
    assign window_rom[371]={1'b0, 13'd6685};
    assign window_rom[372]={1'b0, 13'd6704};
    assign window_rom[373]={1'b0, 13'd6722};
    assign window_rom[374]={1'b0, 13'd6741};
    assign window_rom[375]={1'b0, 13'd6760};
    assign window_rom[376]={1'b0, 13'd6778};
    assign window_rom[377]={1'b0, 13'd6797};
    assign window_rom[378]={1'b0, 13'd6815};
    assign window_rom[379]={1'b0, 13'd6833};
    assign window_rom[380]={1'b0, 13'd6851};
    assign window_rom[381]={1'b0, 13'd6869};
    assign window_rom[382]={1'b0, 13'd6887};
    assign window_rom[383]={1'b0, 13'd6905};
    assign window_rom[384]={1'b0, 13'd6922};
    assign window_rom[385]={1'b0, 13'd6940};
    assign window_rom[386]={1'b0, 13'd6957};
    assign window_rom[387]={1'b0, 13'd6975};
    assign window_rom[388]={1'b0, 13'd6992};
    assign window_rom[389]={1'b0, 13'd7009};
    assign window_rom[390]={1'b0, 13'd7026};
    assign window_rom[391]={1'b0, 13'd7043};
    assign window_rom[392]={1'b0, 13'd7060};
    assign window_rom[393]={1'b0, 13'd7076};
    assign window_rom[394]={1'b0, 13'd7093};
    assign window_rom[395]={1'b0, 13'd7109};
    assign window_rom[396]={1'b0, 13'd7126};
    assign window_rom[397]={1'b0, 13'd7142};
    assign window_rom[398]={1'b0, 13'd7158};
    assign window_rom[399]={1'b0, 13'd7174};
    assign window_rom[400]={1'b0, 13'd7190};
    assign window_rom[401]={1'b0, 13'd7205};
    assign window_rom[402]={1'b0, 13'd7221};
    assign window_rom[403]={1'b0, 13'd7236};
    assign window_rom[404]={1'b0, 13'd7252};
    assign window_rom[405]={1'b0, 13'd7267};
    assign window_rom[406]={1'b0, 13'd7282};
    assign window_rom[407]={1'b0, 13'd7297};
    assign window_rom[408]={1'b0, 13'd7312};
    assign window_rom[409]={1'b0, 13'd7327};
    assign window_rom[410]={1'b0, 13'd7341};
    assign window_rom[411]={1'b0, 13'd7356};
    assign window_rom[412]={1'b0, 13'd7370};
    assign window_rom[413]={1'b0, 13'd7385};
    assign window_rom[414]={1'b0, 13'd7399};
    assign window_rom[415]={1'b0, 13'd7413};
    assign window_rom[416]={1'b0, 13'd7427};
    assign window_rom[417]={1'b0, 13'd7440};
    assign window_rom[418]={1'b0, 13'd7454};
    assign window_rom[419]={1'b0, 13'd7468};
    assign window_rom[420]={1'b0, 13'd7481};
    assign window_rom[421]={1'b0, 13'd7494};
    assign window_rom[422]={1'b0, 13'd7507};
    assign window_rom[423]={1'b0, 13'd7520};
    assign window_rom[424]={1'b0, 13'd7533};
    assign window_rom[425]={1'b0, 13'd7546};
    assign window_rom[426]={1'b0, 13'd7558};
    assign window_rom[427]={1'b0, 13'd7571};
    assign window_rom[428]={1'b0, 13'd7583};
    assign window_rom[429]={1'b0, 13'd7595};
    assign window_rom[430]={1'b0, 13'd7608};
    assign window_rom[431]={1'b0, 13'd7619};
    assign window_rom[432]={1'b0, 13'd7631};
    assign window_rom[433]={1'b0, 13'd7643};
    assign window_rom[434]={1'b0, 13'd7654};
    assign window_rom[435]={1'b0, 13'd7666};
    assign window_rom[436]={1'b0, 13'd7677};
    assign window_rom[437]={1'b0, 13'd7688};
    assign window_rom[438]={1'b0, 13'd7699};
    assign window_rom[439]={1'b0, 13'd7710};
    assign window_rom[440]={1'b0, 13'd7721};
    assign window_rom[441]={1'b0, 13'd7731};
    assign window_rom[442]={1'b0, 13'd7742};
    assign window_rom[443]={1'b0, 13'd7752};
    assign window_rom[444]={1'b0, 13'd7762};
    assign window_rom[445]={1'b0, 13'd7772};
    assign window_rom[446]={1'b0, 13'd7782};
    assign window_rom[447]={1'b0, 13'd7792};
    assign window_rom[448]={1'b0, 13'd7801};
    assign window_rom[449]={1'b0, 13'd7811};
    assign window_rom[450]={1'b0, 13'd7820};
    assign window_rom[451]={1'b0, 13'd7829};
    assign window_rom[452]={1'b0, 13'd7838};
    assign window_rom[453]={1'b0, 13'd7847};
    assign window_rom[454]={1'b0, 13'd7856};
    assign window_rom[455]={1'b0, 13'd7865};
    assign window_rom[456]={1'b0, 13'd7873};
    assign window_rom[457]={1'b0, 13'd7881};
    assign window_rom[458]={1'b0, 13'd7890};
    assign window_rom[459]={1'b0, 13'd7898};
    assign window_rom[460]={1'b0, 13'd7905};
    assign window_rom[461]={1'b0, 13'd7913};
    assign window_rom[462]={1'b0, 13'd7921};
    assign window_rom[463]={1'b0, 13'd7928};
    assign window_rom[464]={1'b0, 13'd7935};
    assign window_rom[465]={1'b0, 13'd7943};
    assign window_rom[466]={1'b0, 13'd7950};
    assign window_rom[467]={1'b0, 13'd7956};
    assign window_rom[468]={1'b0, 13'd7963};
    assign window_rom[469]={1'b0, 13'd7970};
    assign window_rom[470]={1'b0, 13'd7976};
    assign window_rom[471]={1'b0, 13'd7982};
    assign window_rom[472]={1'b0, 13'd7989};
    assign window_rom[473]={1'b0, 13'd7995};
    assign window_rom[474]={1'b0, 13'd8000};
    assign window_rom[475]={1'b0, 13'd8006};
    assign window_rom[476]={1'b0, 13'd8012};
    assign window_rom[477]={1'b0, 13'd8017};
    assign window_rom[478]={1'b0, 13'd8022};
    assign window_rom[479]={1'b0, 13'd8027};
    assign window_rom[480]={1'b0, 13'd8032};
    assign window_rom[481]={1'b0, 13'd8037};
    assign window_rom[482]={1'b0, 13'd8042};
    assign window_rom[483]={1'b0, 13'd8046};
    assign window_rom[484]={1'b0, 13'd8050};
    assign window_rom[485]={1'b0, 13'd8055};
    assign window_rom[486]={1'b0, 13'd8059};
    assign window_rom[487]={1'b0, 13'd8062};
    assign window_rom[488]={1'b0, 13'd8066};
    assign window_rom[489]={1'b0, 13'd8070};
    assign window_rom[490]={1'b0, 13'd8073};
    assign window_rom[491]={1'b0, 13'd8076};
    assign window_rom[492]={1'b0, 13'd8080};
    assign window_rom[493]={1'b0, 13'd8083};
    assign window_rom[494]={1'b0, 13'd8085};
    assign window_rom[495]={1'b0, 13'd8088};
    assign window_rom[496]={1'b0, 13'd8091};
    assign window_rom[497]={1'b0, 13'd8093};
    assign window_rom[498]={1'b0, 13'd8095};
    assign window_rom[499]={1'b0, 13'd8097};
    assign window_rom[500]={1'b0, 13'd8099};
    assign window_rom[501]={1'b0, 13'd8101};
    assign window_rom[502]={1'b0, 13'd8102};
    assign window_rom[503]={1'b0, 13'd8104};
    assign window_rom[504]={1'b0, 13'd8105};
    assign window_rom[505]={1'b0, 13'd8106};
    assign window_rom[506]={1'b0, 13'd8107};
    assign window_rom[507]={1'b0, 13'd8108};
    assign window_rom[508]={1'b0, 13'd8109};
    assign window_rom[509]={1'b0, 13'd8109};
    assign window_rom[510]={1'b0, 13'd8110};
    assign window_rom[511]={1'b0, 13'd8110};
    assign window_rom[512]={1'b0, 13'd8110};
    assign window_rom[513]={1'b0, 13'd8110};
    assign window_rom[514]={1'b0, 13'd8110};
    assign window_rom[515]={1'b0, 13'd8109};
    assign window_rom[516]={1'b0, 13'd8109};
    assign window_rom[517]={1'b0, 13'd8108};
    assign window_rom[518]={1'b0, 13'd8107};
    assign window_rom[519]={1'b0, 13'd8106};
    assign window_rom[520]={1'b0, 13'd8105};
    assign window_rom[521]={1'b0, 13'd8104};
    assign window_rom[522]={1'b0, 13'd8102};
    assign window_rom[523]={1'b0, 13'd8101};
    assign window_rom[524]={1'b0, 13'd8099};
    assign window_rom[525]={1'b0, 13'd8097};
    assign window_rom[526]={1'b0, 13'd8095};
    assign window_rom[527]={1'b0, 13'd8093};
    assign window_rom[528]={1'b0, 13'd8091};
    assign window_rom[529]={1'b0, 13'd8088};
    assign window_rom[530]={1'b0, 13'd8085};
    assign window_rom[531]={1'b0, 13'd8083};
    assign window_rom[532]={1'b0, 13'd8080};
    assign window_rom[533]={1'b0, 13'd8076};
    assign window_rom[534]={1'b0, 13'd8073};
    assign window_rom[535]={1'b0, 13'd8070};
    assign window_rom[536]={1'b0, 13'd8066};
    assign window_rom[537]={1'b0, 13'd8062};
    assign window_rom[538]={1'b0, 13'd8059};
    assign window_rom[539]={1'b0, 13'd8055};
    assign window_rom[540]={1'b0, 13'd8050};
    assign window_rom[541]={1'b0, 13'd8046};
    assign window_rom[542]={1'b0, 13'd8042};
    assign window_rom[543]={1'b0, 13'd8037};
    assign window_rom[544]={1'b0, 13'd8032};
    assign window_rom[545]={1'b0, 13'd8027};
    assign window_rom[546]={1'b0, 13'd8022};
    assign window_rom[547]={1'b0, 13'd8017};
    assign window_rom[548]={1'b0, 13'd8012};
    assign window_rom[549]={1'b0, 13'd8006};
    assign window_rom[550]={1'b0, 13'd8000};
    assign window_rom[551]={1'b0, 13'd7995};
    assign window_rom[552]={1'b0, 13'd7989};
    assign window_rom[553]={1'b0, 13'd7982};
    assign window_rom[554]={1'b0, 13'd7976};
    assign window_rom[555]={1'b0, 13'd7970};
    assign window_rom[556]={1'b0, 13'd7963};
    assign window_rom[557]={1'b0, 13'd7956};
    assign window_rom[558]={1'b0, 13'd7950};
    assign window_rom[559]={1'b0, 13'd7943};
    assign window_rom[560]={1'b0, 13'd7935};
    assign window_rom[561]={1'b0, 13'd7928};
    assign window_rom[562]={1'b0, 13'd7921};
    assign window_rom[563]={1'b0, 13'd7913};
    assign window_rom[564]={1'b0, 13'd7905};
    assign window_rom[565]={1'b0, 13'd7898};
    assign window_rom[566]={1'b0, 13'd7890};
    assign window_rom[567]={1'b0, 13'd7881};
    assign window_rom[568]={1'b0, 13'd7873};
    assign window_rom[569]={1'b0, 13'd7865};
    assign window_rom[570]={1'b0, 13'd7856};
    assign window_rom[571]={1'b0, 13'd7847};
    assign window_rom[572]={1'b0, 13'd7838};
    assign window_rom[573]={1'b0, 13'd7829};
    assign window_rom[574]={1'b0, 13'd7820};
    assign window_rom[575]={1'b0, 13'd7811};
    assign window_rom[576]={1'b0, 13'd7801};
    assign window_rom[577]={1'b0, 13'd7792};
    assign window_rom[578]={1'b0, 13'd7782};
    assign window_rom[579]={1'b0, 13'd7772};
    assign window_rom[580]={1'b0, 13'd7762};
    assign window_rom[581]={1'b0, 13'd7752};
    assign window_rom[582]={1'b0, 13'd7742};
    assign window_rom[583]={1'b0, 13'd7731};
    assign window_rom[584]={1'b0, 13'd7721};
    assign window_rom[585]={1'b0, 13'd7710};
    assign window_rom[586]={1'b0, 13'd7699};
    assign window_rom[587]={1'b0, 13'd7688};
    assign window_rom[588]={1'b0, 13'd7677};
    assign window_rom[589]={1'b0, 13'd7666};
    assign window_rom[590]={1'b0, 13'd7654};
    assign window_rom[591]={1'b0, 13'd7643};
    assign window_rom[592]={1'b0, 13'd7631};
    assign window_rom[593]={1'b0, 13'd7619};
    assign window_rom[594]={1'b0, 13'd7608};
    assign window_rom[595]={1'b0, 13'd7595};
    assign window_rom[596]={1'b0, 13'd7583};
    assign window_rom[597]={1'b0, 13'd7571};
    assign window_rom[598]={1'b0, 13'd7558};
    assign window_rom[599]={1'b0, 13'd7546};
    assign window_rom[600]={1'b0, 13'd7533};
    assign window_rom[601]={1'b0, 13'd7520};
    assign window_rom[602]={1'b0, 13'd7507};
    assign window_rom[603]={1'b0, 13'd7494};
    assign window_rom[604]={1'b0, 13'd7481};
    assign window_rom[605]={1'b0, 13'd7468};
    assign window_rom[606]={1'b0, 13'd7454};
    assign window_rom[607]={1'b0, 13'd7440};
    assign window_rom[608]={1'b0, 13'd7427};
    assign window_rom[609]={1'b0, 13'd7413};
    assign window_rom[610]={1'b0, 13'd7399};
    assign window_rom[611]={1'b0, 13'd7385};
    assign window_rom[612]={1'b0, 13'd7370};
    assign window_rom[613]={1'b0, 13'd7356};
    assign window_rom[614]={1'b0, 13'd7341};
    assign window_rom[615]={1'b0, 13'd7327};
    assign window_rom[616]={1'b0, 13'd7312};
    assign window_rom[617]={1'b0, 13'd7297};
    assign window_rom[618]={1'b0, 13'd7282};
    assign window_rom[619]={1'b0, 13'd7267};
    assign window_rom[620]={1'b0, 13'd7252};
    assign window_rom[621]={1'b0, 13'd7236};
    assign window_rom[622]={1'b0, 13'd7221};
    assign window_rom[623]={1'b0, 13'd7205};
    assign window_rom[624]={1'b0, 13'd7190};
    assign window_rom[625]={1'b0, 13'd7174};
    assign window_rom[626]={1'b0, 13'd7158};
    assign window_rom[627]={1'b0, 13'd7142};
    assign window_rom[628]={1'b0, 13'd7126};
    assign window_rom[629]={1'b0, 13'd7109};
    assign window_rom[630]={1'b0, 13'd7093};
    assign window_rom[631]={1'b0, 13'd7076};
    assign window_rom[632]={1'b0, 13'd7060};
    assign window_rom[633]={1'b0, 13'd7043};
    assign window_rom[634]={1'b0, 13'd7026};
    assign window_rom[635]={1'b0, 13'd7009};
    assign window_rom[636]={1'b0, 13'd6992};
    assign window_rom[637]={1'b0, 13'd6975};
    assign window_rom[638]={1'b0, 13'd6957};
    assign window_rom[639]={1'b0, 13'd6940};
    assign window_rom[640]={1'b0, 13'd6922};
    assign window_rom[641]={1'b0, 13'd6905};
    assign window_rom[642]={1'b0, 13'd6887};
    assign window_rom[643]={1'b0, 13'd6869};
    assign window_rom[644]={1'b0, 13'd6851};
    assign window_rom[645]={1'b0, 13'd6833};
    assign window_rom[646]={1'b0, 13'd6815};
    assign window_rom[647]={1'b0, 13'd6797};
    assign window_rom[648]={1'b0, 13'd6778};
    assign window_rom[649]={1'b0, 13'd6760};
    assign window_rom[650]={1'b0, 13'd6741};
    assign window_rom[651]={1'b0, 13'd6722};
    assign window_rom[652]={1'b0, 13'd6704};
    assign window_rom[653]={1'b0, 13'd6685};
    assign window_rom[654]={1'b0, 13'd6666};
    assign window_rom[655]={1'b0, 13'd6647};
    assign window_rom[656]={1'b0, 13'd6628};
    assign window_rom[657]={1'b0, 13'd6608};
    assign window_rom[658]={1'b0, 13'd6589};
    assign window_rom[659]={1'b0, 13'd6569};
    assign window_rom[660]={1'b0, 13'd6550};
    assign window_rom[661]={1'b0, 13'd6530};
    assign window_rom[662]={1'b0, 13'd6510};
    assign window_rom[663]={1'b0, 13'd6491};
    assign window_rom[664]={1'b0, 13'd6471};
    assign window_rom[665]={1'b0, 13'd6451};
    assign window_rom[666]={1'b0, 13'd6430};
    assign window_rom[667]={1'b0, 13'd6410};
    assign window_rom[668]={1'b0, 13'd6390};
    assign window_rom[669]={1'b0, 13'd6370};
    assign window_rom[670]={1'b0, 13'd6349};
    assign window_rom[671]={1'b0, 13'd6329};
    assign window_rom[672]={1'b0, 13'd6308};
    assign window_rom[673]={1'b0, 13'd6287};
    assign window_rom[674]={1'b0, 13'd6266};
    assign window_rom[675]={1'b0, 13'd6245};
    assign window_rom[676]={1'b0, 13'd6224};
    assign window_rom[677]={1'b0, 13'd6203};
    assign window_rom[678]={1'b0, 13'd6182};
    assign window_rom[679]={1'b0, 13'd6161};
    assign window_rom[680]={1'b0, 13'd6140};
    assign window_rom[681]={1'b0, 13'd6118};
    assign window_rom[682]={1'b0, 13'd6097};
    assign window_rom[683]={1'b0, 13'd6075};
    assign window_rom[684]={1'b0, 13'd6054};
    assign window_rom[685]={1'b0, 13'd6032};
    assign window_rom[686]={1'b0, 13'd6010};
    assign window_rom[687]={1'b0, 13'd5988};
    assign window_rom[688]={1'b0, 13'd5967};
    assign window_rom[689]={1'b0, 13'd5945};
    assign window_rom[690]={1'b0, 13'd5923};
    assign window_rom[691]={1'b0, 13'd5900};
    assign window_rom[692]={1'b0, 13'd5878};
    assign window_rom[693]={1'b0, 13'd5856};
    assign window_rom[694]={1'b0, 13'd5834};
    assign window_rom[695]={1'b0, 13'd5811};
    assign window_rom[696]={1'b0, 13'd5789};
    assign window_rom[697]={1'b0, 13'd5766};
    assign window_rom[698]={1'b0, 13'd5744};
    assign window_rom[699]={1'b0, 13'd5721};
    assign window_rom[700]={1'b0, 13'd5698};
    assign window_rom[701]={1'b0, 13'd5676};
    assign window_rom[702]={1'b0, 13'd5653};
    assign window_rom[703]={1'b0, 13'd5630};
    assign window_rom[704]={1'b0, 13'd5607};
    assign window_rom[705]={1'b0, 13'd5584};
    assign window_rom[706]={1'b0, 13'd5561};
    assign window_rom[707]={1'b0, 13'd5538};
    assign window_rom[708]={1'b0, 13'd5514};
    assign window_rom[709]={1'b0, 13'd5491};
    assign window_rom[710]={1'b0, 13'd5468};
    assign window_rom[711]={1'b0, 13'd5445};
    assign window_rom[712]={1'b0, 13'd5421};
    assign window_rom[713]={1'b0, 13'd5398};
    assign window_rom[714]={1'b0, 13'd5374};
    assign window_rom[715]={1'b0, 13'd5351};
    assign window_rom[716]={1'b0, 13'd5327};
    assign window_rom[717]={1'b0, 13'd5303};
    assign window_rom[718]={1'b0, 13'd5280};
    assign window_rom[719]={1'b0, 13'd5256};
    assign window_rom[720]={1'b0, 13'd5232};
    assign window_rom[721]={1'b0, 13'd5208};
    assign window_rom[722]={1'b0, 13'd5184};
    assign window_rom[723]={1'b0, 13'd5161};
    assign window_rom[724]={1'b0, 13'd5137};
    assign window_rom[725]={1'b0, 13'd5113};
    assign window_rom[726]={1'b0, 13'd5089};
    assign window_rom[727]={1'b0, 13'd5064};
    assign window_rom[728]={1'b0, 13'd5040};
    assign window_rom[729]={1'b0, 13'd5016};
    assign window_rom[730]={1'b0, 13'd4992};
    assign window_rom[731]={1'b0, 13'd4968};
    assign window_rom[732]={1'b0, 13'd4944};
    assign window_rom[733]={1'b0, 13'd4919};
    assign window_rom[734]={1'b0, 13'd4895};
    assign window_rom[735]={1'b0, 13'd4871};
    assign window_rom[736]={1'b0, 13'd4846};
    assign window_rom[737]={1'b0, 13'd4822};
    assign window_rom[738]={1'b0, 13'd4797};
    assign window_rom[739]={1'b0, 13'd4773};
    assign window_rom[740]={1'b0, 13'd4748};
    assign window_rom[741]={1'b0, 13'd4724};
    assign window_rom[742]={1'b0, 13'd4699};
    assign window_rom[743]={1'b0, 13'd4675};
    assign window_rom[744]={1'b0, 13'd4650};
    assign window_rom[745]={1'b0, 13'd4625};
    assign window_rom[746]={1'b0, 13'd4601};
    assign window_rom[747]={1'b0, 13'd4576};
    assign window_rom[748]={1'b0, 13'd4551};
    assign window_rom[749]={1'b0, 13'd4527};
    assign window_rom[750]={1'b0, 13'd4502};
    assign window_rom[751]={1'b0, 13'd4477};
    assign window_rom[752]={1'b0, 13'd4453};
    assign window_rom[753]={1'b0, 13'd4428};
    assign window_rom[754]={1'b0, 13'd4403};
    assign window_rom[755]={1'b0, 13'd4378};
    assign window_rom[756]={1'b0, 13'd4353};
    assign window_rom[757]={1'b0, 13'd4329};
    assign window_rom[758]={1'b0, 13'd4304};
    assign window_rom[759]={1'b0, 13'd4279};
    assign window_rom[760]={1'b0, 13'd4254};
    assign window_rom[761]={1'b0, 13'd4229};
    assign window_rom[762]={1'b0, 13'd4204};
    assign window_rom[763]={1'b0, 13'd4179};
    assign window_rom[764]={1'b0, 13'd4155};
    assign window_rom[765]={1'b0, 13'd4130};
    assign window_rom[766]={1'b0, 13'd4105};
    assign window_rom[767]={1'b0, 13'd4080};
    assign window_rom[768]={1'b0, 13'd4055};
    assign window_rom[769]={1'b0, 13'd4030};
    assign window_rom[770]={1'b0, 13'd4005};
    assign window_rom[771]={1'b0, 13'd3980};
    assign window_rom[772]={1'b0, 13'd3956};
    assign window_rom[773]={1'b0, 13'd3931};
    assign window_rom[774]={1'b0, 13'd3906};
    assign window_rom[775]={1'b0, 13'd3881};
    assign window_rom[776]={1'b0, 13'd3856};
    assign window_rom[777]={1'b0, 13'd3831};
    assign window_rom[778]={1'b0, 13'd3806};
    assign window_rom[779]={1'b0, 13'd3782};
    assign window_rom[780]={1'b0, 13'd3757};
    assign window_rom[781]={1'b0, 13'd3732};
    assign window_rom[782]={1'b0, 13'd3707};
    assign window_rom[783]={1'b0, 13'd3682};
    assign window_rom[784]={1'b0, 13'd3658};
    assign window_rom[785]={1'b0, 13'd3633};
    assign window_rom[786]={1'b0, 13'd3608};
    assign window_rom[787]={1'b0, 13'd3583};
    assign window_rom[788]={1'b0, 13'd3559};
    assign window_rom[789]={1'b0, 13'd3534};
    assign window_rom[790]={1'b0, 13'd3509};
    assign window_rom[791]={1'b0, 13'd3485};
    assign window_rom[792]={1'b0, 13'd3460};
    assign window_rom[793]={1'b0, 13'd3435};
    assign window_rom[794]={1'b0, 13'd3411};
    assign window_rom[795]={1'b0, 13'd3386};
    assign window_rom[796]={1'b0, 13'd3362};
    assign window_rom[797]={1'b0, 13'd3337};
    assign window_rom[798]={1'b0, 13'd3313};
    assign window_rom[799]={1'b0, 13'd3288};
    assign window_rom[800]={1'b0, 13'd3264};
    assign window_rom[801]={1'b0, 13'd3240};
    assign window_rom[802]={1'b0, 13'd3215};
    assign window_rom[803]={1'b0, 13'd3191};
    assign window_rom[804]={1'b0, 13'd3167};
    assign window_rom[805]={1'b0, 13'd3142};
    assign window_rom[806]={1'b0, 13'd3118};
    assign window_rom[807]={1'b0, 13'd3094};
    assign window_rom[808]={1'b0, 13'd3070};
    assign window_rom[809]={1'b0, 13'd3046};
    assign window_rom[810]={1'b0, 13'd3022};
    assign window_rom[811]={1'b0, 13'd2998};
    assign window_rom[812]={1'b0, 13'd2974};
    assign window_rom[813]={1'b0, 13'd2950};
    assign window_rom[814]={1'b0, 13'd2926};
    assign window_rom[815]={1'b0, 13'd2902};
    assign window_rom[816]={1'b0, 13'd2878};
    assign window_rom[817]={1'b0, 13'd2854};
    assign window_rom[818]={1'b0, 13'd2830};
    assign window_rom[819]={1'b0, 13'd2807};
    assign window_rom[820]={1'b0, 13'd2783};
    assign window_rom[821]={1'b0, 13'd2759};
    assign window_rom[822]={1'b0, 13'd2736};
    assign window_rom[823]={1'b0, 13'd2712};
    assign window_rom[824]={1'b0, 13'd2689};
    assign window_rom[825]={1'b0, 13'd2666};
    assign window_rom[826]={1'b0, 13'd2642};
    assign window_rom[827]={1'b0, 13'd2619};
    assign window_rom[828]={1'b0, 13'd2596};
    assign window_rom[829]={1'b0, 13'd2572};
    assign window_rom[830]={1'b0, 13'd2549};
    assign window_rom[831]={1'b0, 13'd2526};
    assign window_rom[832]={1'b0, 13'd2503};
    assign window_rom[833]={1'b0, 13'd2480};
    assign window_rom[834]={1'b0, 13'd2457};
    assign window_rom[835]={1'b0, 13'd2435};
    assign window_rom[836]={1'b0, 13'd2412};
    assign window_rom[837]={1'b0, 13'd2389};
    assign window_rom[838]={1'b0, 13'd2366};
    assign window_rom[839]={1'b0, 13'd2344};
    assign window_rom[840]={1'b0, 13'd2321};
    assign window_rom[841]={1'b0, 13'd2299};
    assign window_rom[842]={1'b0, 13'd2276};
    assign window_rom[843]={1'b0, 13'd2254};
    assign window_rom[844]={1'b0, 13'd2232};
    assign window_rom[845]={1'b0, 13'd2210};
    assign window_rom[846]={1'b0, 13'd2188};
    assign window_rom[847]={1'b0, 13'd2165};
    assign window_rom[848]={1'b0, 13'd2144};
    assign window_rom[849]={1'b0, 13'd2122};
    assign window_rom[850]={1'b0, 13'd2100};
    assign window_rom[851]={1'b0, 13'd2078};
    assign window_rom[852]={1'b0, 13'd2056};
    assign window_rom[853]={1'b0, 13'd2035};
    assign window_rom[854]={1'b0, 13'd2013};
    assign window_rom[855]={1'b0, 13'd1992};
    assign window_rom[856]={1'b0, 13'd1970};
    assign window_rom[857]={1'b0, 13'd1949};
    assign window_rom[858]={1'b0, 13'd1928};
    assign window_rom[859]={1'b0, 13'd1907};
    assign window_rom[860]={1'b0, 13'd1886};
    assign window_rom[861]={1'b0, 13'd1865};
    assign window_rom[862]={1'b0, 13'd1844};
    assign window_rom[863]={1'b0, 13'd1823};
    assign window_rom[864]={1'b0, 13'd1802};
    assign window_rom[865]={1'b0, 13'd1782};
    assign window_rom[866]={1'b0, 13'd1761};
    assign window_rom[867]={1'b0, 13'd1741};
    assign window_rom[868]={1'b0, 13'd1720};
    assign window_rom[869]={1'b0, 13'd1700};
    assign window_rom[870]={1'b0, 13'd1680};
    assign window_rom[871]={1'b0, 13'd1659};
    assign window_rom[872]={1'b0, 13'd1639};
    assign window_rom[873]={1'b0, 13'd1620};
    assign window_rom[874]={1'b0, 13'd1600};
    assign window_rom[875]={1'b0, 13'd1580};
    assign window_rom[876]={1'b0, 13'd1560};
    assign window_rom[877]={1'b0, 13'd1541};
    assign window_rom[878]={1'b0, 13'd1521};
    assign window_rom[879]={1'b0, 13'd1502};
    assign window_rom[880]={1'b0, 13'd1483};
    assign window_rom[881]={1'b0, 13'd1463};
    assign window_rom[882]={1'b0, 13'd1444};
    assign window_rom[883]={1'b0, 13'd1425};
    assign window_rom[884]={1'b0, 13'd1406};
    assign window_rom[885]={1'b0, 13'd1388};
    assign window_rom[886]={1'b0, 13'd1369};
    assign window_rom[887]={1'b0, 13'd1350};
    assign window_rom[888]={1'b0, 13'd1332};
    assign window_rom[889]={1'b0, 13'd1313};
    assign window_rom[890]={1'b0, 13'd1295};
    assign window_rom[891]={1'b0, 13'd1277};
    assign window_rom[892]={1'b0, 13'd1259};
    assign window_rom[893]={1'b0, 13'd1241};
    assign window_rom[894]={1'b0, 13'd1223};
    assign window_rom[895]={1'b0, 13'd1205};
    assign window_rom[896]={1'b0, 13'd1188};
    assign window_rom[897]={1'b0, 13'd1170};
    assign window_rom[898]={1'b0, 13'd1153};
    assign window_rom[899]={1'b0, 13'd1135};
    assign window_rom[900]={1'b0, 13'd1118};
    assign window_rom[901]={1'b0, 13'd1101};
    assign window_rom[902]={1'b0, 13'd1084};
    assign window_rom[903]={1'b0, 13'd1067};
    assign window_rom[904]={1'b0, 13'd1050};
    assign window_rom[905]={1'b0, 13'd1034};
    assign window_rom[906]={1'b0, 13'd1017};
    assign window_rom[907]={1'b0, 13'd1001};
    assign window_rom[908]={1'b0, 13'd985};
    assign window_rom[909]={1'b0, 13'd968};
    assign window_rom[910]={1'b0, 13'd952};
    assign window_rom[911]={1'b0, 13'd936};
    assign window_rom[912]={1'b0, 13'd920};
    assign window_rom[913]={1'b0, 13'd905};
    assign window_rom[914]={1'b0, 13'd889};
    assign window_rom[915]={1'b0, 13'd874};
    assign window_rom[916]={1'b0, 13'd858};
    assign window_rom[917]={1'b0, 13'd843};
    assign window_rom[918]={1'b0, 13'd828};
    assign window_rom[919]={1'b0, 13'd813};
    assign window_rom[920]={1'b0, 13'd798};
    assign window_rom[921]={1'b0, 13'd783};
    assign window_rom[922]={1'b0, 13'd769};
    assign window_rom[923]={1'b0, 13'd754};
    assign window_rom[924]={1'b0, 13'd740};
    assign window_rom[925]={1'b0, 13'd725};
    assign window_rom[926]={1'b0, 13'd711};
    assign window_rom[927]={1'b0, 13'd697};
    assign window_rom[928]={1'b0, 13'd683};
    assign window_rom[929]={1'b0, 13'd670};
    assign window_rom[930]={1'b0, 13'd656};
    assign window_rom[931]={1'b0, 13'd643};
    assign window_rom[932]={1'b0, 13'd629};
    assign window_rom[933]={1'b0, 13'd616};
    assign window_rom[934]={1'b0, 13'd603};
    assign window_rom[935]={1'b0, 13'd590};
    assign window_rom[936]={1'b0, 13'd577};
    assign window_rom[937]={1'b0, 13'd564};
    assign window_rom[938]={1'b0, 13'd552};
    assign window_rom[939]={1'b0, 13'd539};
    assign window_rom[940]={1'b0, 13'd527};
    assign window_rom[941]={1'b0, 13'd515};
    assign window_rom[942]={1'b0, 13'd503};
    assign window_rom[943]={1'b0, 13'd491};
    assign window_rom[944]={1'b0, 13'd479};
    assign window_rom[945]={1'b0, 13'd467};
    assign window_rom[946]={1'b0, 13'd456};
    assign window_rom[947]={1'b0, 13'd444};
    assign window_rom[948]={1'b0, 13'd433};
    assign window_rom[949]={1'b0, 13'd422};
    assign window_rom[950]={1'b0, 13'd411};
    assign window_rom[951]={1'b0, 13'd400};
    assign window_rom[952]={1'b0, 13'd389};
    assign window_rom[953]={1'b0, 13'd379};
    assign window_rom[954]={1'b0, 13'd368};
    assign window_rom[955]={1'b0, 13'd358};
    assign window_rom[956]={1'b0, 13'd348};
    assign window_rom[957]={1'b0, 13'd338};
    assign window_rom[958]={1'b0, 13'd328};
    assign window_rom[959]={1'b0, 13'd318};
    assign window_rom[960]={1'b0, 13'd309};
    assign window_rom[961]={1'b0, 13'd299};
    assign window_rom[962]={1'b0, 13'd290};
    assign window_rom[963]={1'b0, 13'd281};
    assign window_rom[964]={1'b0, 13'd272};
    assign window_rom[965]={1'b0, 13'd263};
    assign window_rom[966]={1'b0, 13'd254};
    assign window_rom[967]={1'b0, 13'd245};
    assign window_rom[968]={1'b0, 13'd237};
    assign window_rom[969]={1'b0, 13'd229};
    assign window_rom[970]={1'b0, 13'd221};
    assign window_rom[971]={1'b0, 13'd213};
    assign window_rom[972]={1'b0, 13'd205};
    assign window_rom[973]={1'b0, 13'd197};
    assign window_rom[974]={1'b0, 13'd189};
    assign window_rom[975]={1'b0, 13'd182};
    assign window_rom[976]={1'b0, 13'd175};
    assign window_rom[977]={1'b0, 13'd167};
    assign window_rom[978]={1'b0, 13'd160};
    assign window_rom[979]={1'b0, 13'd154};
    assign window_rom[980]={1'b0, 13'd147};
    assign window_rom[981]={1'b0, 13'd140};
    assign window_rom[982]={1'b0, 13'd134};
    assign window_rom[983]={1'b0, 13'd128};
    assign window_rom[984]={1'b0, 13'd122};
    assign window_rom[985]={1'b0, 13'd116};
    assign window_rom[986]={1'b0, 13'd110};
    assign window_rom[987]={1'b0, 13'd104};
    assign window_rom[988]={1'b0, 13'd99};
    assign window_rom[989]={1'b0, 13'd93};
    assign window_rom[990]={1'b0, 13'd88};
    assign window_rom[991]={1'b0, 13'd83};
    assign window_rom[992]={1'b0, 13'd78};
    assign window_rom[993]={1'b0, 13'd73};
    assign window_rom[994]={1'b0, 13'd69};
    assign window_rom[995]={1'b0, 13'd64};
    assign window_rom[996]={1'b0, 13'd60};
    assign window_rom[997]={1'b0, 13'd56};
    assign window_rom[998]={1'b0, 13'd51};
    assign window_rom[999]={1'b0, 13'd48};
    assign window_rom[1000]={1'b0, 13'd44};
    assign window_rom[1001]={1'b0, 13'd40};
    assign window_rom[1002]={1'b0, 13'd37};
    assign window_rom[1003]={1'b0, 13'd34};
    assign window_rom[1004]={1'b0, 13'd30};
    assign window_rom[1005]={1'b0, 13'd28};
    assign window_rom[1006]={1'b0, 13'd25};
    assign window_rom[1007]={1'b0, 13'd22};
    assign window_rom[1008]={1'b0, 13'd20};
    assign window_rom[1009]={1'b0, 13'd17};
    assign window_rom[1010]={1'b0, 13'd15};
    assign window_rom[1011]={1'b0, 13'd13};
    assign window_rom[1012]={1'b0, 13'd11};
    assign window_rom[1013]={1'b0, 13'd9};
    assign window_rom[1014]={1'b0, 13'd8};
    assign window_rom[1015]={1'b0, 13'd6};
    assign window_rom[1016]={1'b0, 13'd5};
    assign window_rom[1017]={1'b0, 13'd4};
    assign window_rom[1018]={1'b0, 13'd3};
    assign window_rom[1019]={1'b0, 13'd2};
    assign window_rom[1020]={1'b0, 13'd1};
    assign window_rom[1021]={1'b0, 13'd1};
    assign window_rom[1022]={1'b0, 13'd0};
    assign window_rom[1023]={1'b0, 13'd0};

endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */