module mel_rom (
    input  wire               clk,
    input  wire               rst_n,
    input  wire        [ 9:0] addr,
    input  wire               in_nd,
    output reg signed [ 39:0] w
  );

reg [39:0] dout [0:1023];


initial begin
dout[0]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[1]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[2]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[3]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[4]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[5]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[6]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[7]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[8]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[9]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[10]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[11]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[12]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[13]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[14]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[15]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[16]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[17]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[18]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[19]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[20]={ 4'd1     ,  4'd0, 16'd4681   ,16'd0};
dout[21]={ 4'd1     ,  4'd0, 16'd9362   ,16'd0};
dout[22]={ 4'd1     ,  4'd0, 16'd14043   ,16'd0};
dout[23]={ 4'd1     ,  4'd0, 16'd18724   ,16'd0};
dout[24]={ 4'd1     ,  4'd0, 16'd23405   ,16'd0};
dout[25]={ 4'd1     ,  4'd0, 16'd28086   ,16'd0};
dout[26]={ 4'd1     ,  4'd0, 16'd32768   ,16'd0};
dout[27]={ 4'd1     ,  4'd0, 16'd37449   ,16'd0};
dout[28]={ 4'd1     ,  4'd0, 16'd42130   ,16'd0};
dout[29]={ 4'd1     ,  4'd0, 16'd46811   ,16'd0};
dout[30]={ 4'd1     ,  4'd0, 16'd51492   ,16'd0};
dout[31]={ 4'd1     ,  4'd0, 16'd56173   ,16'd0};
dout[32]={ 4'd1     ,  4'd0, 16'd60854   ,16'd0};
dout[33]={ 4'd1     ,  4'd0, 16'd65535   ,16'd0};
dout[34]={ 4'd1     ,  4'd2, 16'd61680   ,16'd3855};
dout[35]={ 4'd1     ,  4'd2, 16'd57825   ,16'd7710};
dout[36]={ 4'd1     ,  4'd2, 16'd53970   ,16'd11565};
dout[37]={ 4'd1     ,  4'd2, 16'd50115   ,16'd15420};
dout[38]={ 4'd1     ,  4'd2, 16'd46260   ,16'd19275};
dout[39]={ 4'd1     ,  4'd2, 16'd42405   ,16'd23130};
dout[40]={ 4'd1     ,  4'd2, 16'd38550   ,16'd26985};
dout[41]={ 4'd1     ,  4'd2, 16'd34695   ,16'd30840};
dout[42]={ 4'd1     ,  4'd2, 16'd30840   ,16'd34695};
dout[43]={ 4'd1     ,  4'd2, 16'd26985   ,16'd38550};
dout[44]={ 4'd1     ,  4'd2, 16'd23130   ,16'd42405};
dout[45]={ 4'd1     ,  4'd2, 16'd19275   ,16'd46260};
dout[46]={ 4'd1     ,  4'd2, 16'd15420   ,16'd50115};
dout[47]={ 4'd1     ,  4'd2, 16'd11565   ,16'd53970};
dout[48]={ 4'd1     ,  4'd2, 16'd7710   ,16'd57825};
dout[49]={ 4'd1     ,  4'd2, 16'd3855   ,16'd61680};
dout[50]={ 4'd2     ,  4'd0, 16'd65535   ,16'd0};
dout[51]={ 4'd2     ,  4'd3, 16'd62259   ,16'd3276};
dout[52]={ 4'd2     ,  4'd3, 16'd58982   ,16'd6553};
dout[53]={ 4'd2     ,  4'd3, 16'd55705   ,16'd9830};
dout[54]={ 4'd2     ,  4'd3, 16'd52428   ,16'd13107};
dout[55]={ 4'd2     ,  4'd3, 16'd49152   ,16'd16384};
dout[56]={ 4'd2     ,  4'd3, 16'd45875   ,16'd19660};
dout[57]={ 4'd2     ,  4'd3, 16'd42598   ,16'd22937};
dout[58]={ 4'd2     ,  4'd3, 16'd39321   ,16'd26214};
dout[59]={ 4'd2     ,  4'd3, 16'd36044   ,16'd29491};
dout[60]={ 4'd2     ,  4'd3, 16'd32768   ,16'd32768};
dout[61]={ 4'd2     ,  4'd3, 16'd29491   ,16'd36044};
dout[62]={ 4'd2     ,  4'd3, 16'd26214   ,16'd39321};
dout[63]={ 4'd2     ,  4'd3, 16'd22937   ,16'd42598};
dout[64]={ 4'd2     ,  4'd3, 16'd19660   ,16'd45875};
dout[65]={ 4'd2     ,  4'd3, 16'd16384   ,16'd49152};
dout[66]={ 4'd2     ,  4'd3, 16'd13107   ,16'd52428};
dout[67]={ 4'd2     ,  4'd3, 16'd9830   ,16'd55705};
dout[68]={ 4'd2     ,  4'd3, 16'd6553   ,16'd58982};
dout[69]={ 4'd2     ,  4'd3, 16'd3276   ,16'd62259};
dout[70]={ 4'd3     ,  4'd0, 16'd65535   ,16'd0};
dout[71]={ 4'd3     ,  4'd4, 16'd62914   ,16'd2621};
dout[72]={ 4'd3     ,  4'd4, 16'd60293   ,16'd5242};
dout[73]={ 4'd3     ,  4'd4, 16'd57671   ,16'd7864};
dout[74]={ 4'd3     ,  4'd4, 16'd55050   ,16'd10485};
dout[75]={ 4'd3     ,  4'd4, 16'd52428   ,16'd13107};
dout[76]={ 4'd3     ,  4'd4, 16'd49807   ,16'd15728};
dout[77]={ 4'd3     ,  4'd4, 16'd47185   ,16'd18350};
dout[78]={ 4'd3     ,  4'd4, 16'd44564   ,16'd20971};
dout[79]={ 4'd3     ,  4'd4, 16'd41943   ,16'd23592};
dout[80]={ 4'd3     ,  4'd4, 16'd39321   ,16'd26214};
dout[81]={ 4'd3     ,  4'd4, 16'd36700   ,16'd28835};
dout[82]={ 4'd3     ,  4'd4, 16'd34078   ,16'd31457};
dout[83]={ 4'd3     ,  4'd4, 16'd31457   ,16'd34078};
dout[84]={ 4'd3     ,  4'd4, 16'd28835   ,16'd36700};
dout[85]={ 4'd3     ,  4'd4, 16'd26214   ,16'd39321};
dout[86]={ 4'd3     ,  4'd4, 16'd23592   ,16'd41943};
dout[87]={ 4'd3     ,  4'd4, 16'd20971   ,16'd44564};
dout[88]={ 4'd3     ,  4'd4, 16'd18350   ,16'd47185};
dout[89]={ 4'd3     ,  4'd4, 16'd15728   ,16'd49807};
dout[90]={ 4'd3     ,  4'd4, 16'd13107   ,16'd52428};
dout[91]={ 4'd3     ,  4'd4, 16'd10485   ,16'd55050};
dout[92]={ 4'd3     ,  4'd4, 16'd7864   ,16'd57671};
dout[93]={ 4'd3     ,  4'd4, 16'd5242   ,16'd60293};
dout[94]={ 4'd3     ,  4'd4, 16'd2621   ,16'd62914};
dout[95]={ 4'd4     ,  4'd0, 16'd65535   ,16'd0};
dout[96]={ 4'd4     ,  4'd5, 16'd63421   ,16'd2114};
dout[97]={ 4'd4     ,  4'd5, 16'd61307   ,16'd4228};
dout[98]={ 4'd4     ,  4'd5, 16'd59193   ,16'd6342};
dout[99]={ 4'd4     ,  4'd5, 16'd57079   ,16'd8456};
dout[100]={ 4'd4     ,  4'd5, 16'd54965   ,16'd10570};
dout[101]={ 4'd4     ,  4'd5, 16'd52851   ,16'd12684};
dout[102]={ 4'd4     ,  4'd5, 16'd50737   ,16'd14798};
dout[103]={ 4'd4     ,  4'd5, 16'd48623   ,16'd16912};
dout[104]={ 4'd4     ,  4'd5, 16'd46509   ,16'd19026};
dout[105]={ 4'd4     ,  4'd5, 16'd44395   ,16'd21140};
dout[106]={ 4'd4     ,  4'd5, 16'd42281   ,16'd23254};
dout[107]={ 4'd4     ,  4'd5, 16'd40167   ,16'd25368};
dout[108]={ 4'd4     ,  4'd5, 16'd38053   ,16'd27482};
dout[109]={ 4'd4     ,  4'd5, 16'd35939   ,16'd29596};
dout[110]={ 4'd4     ,  4'd5, 16'd33825   ,16'd31710};
dout[111]={ 4'd4     ,  4'd5, 16'd31710   ,16'd33825};
dout[112]={ 4'd4     ,  4'd5, 16'd29596   ,16'd35939};
dout[113]={ 4'd4     ,  4'd5, 16'd27482   ,16'd38053};
dout[114]={ 4'd4     ,  4'd5, 16'd25368   ,16'd40167};
dout[115]={ 4'd4     ,  4'd5, 16'd23254   ,16'd42281};
dout[116]={ 4'd4     ,  4'd5, 16'd21140   ,16'd44395};
dout[117]={ 4'd4     ,  4'd5, 16'd19026   ,16'd46509};
dout[118]={ 4'd4     ,  4'd5, 16'd16912   ,16'd48623};
dout[119]={ 4'd4     ,  4'd5, 16'd14798   ,16'd50737};
dout[120]={ 4'd4     ,  4'd5, 16'd12684   ,16'd52851};
dout[121]={ 4'd4     ,  4'd5, 16'd10570   ,16'd54965};
dout[122]={ 4'd4     ,  4'd5, 16'd8456   ,16'd57079};
dout[123]={ 4'd4     ,  4'd5, 16'd6342   ,16'd59193};
dout[124]={ 4'd4     ,  4'd5, 16'd4228   ,16'd61307};
dout[125]={ 4'd4     ,  4'd5, 16'd2114   ,16'd63421};
dout[126]={ 4'd5     ,  4'd0, 16'd65535   ,16'd0};
dout[127]={ 4'd5     ,  4'd6, 16'd63764   ,16'd1771};
dout[128]={ 4'd5     ,  4'd6, 16'd61993   ,16'd3542};
dout[129]={ 4'd5     ,  4'd6, 16'd60222   ,16'd5313};
dout[130]={ 4'd5     ,  4'd6, 16'd58451   ,16'd7084};
dout[131]={ 4'd5     ,  4'd6, 16'd56679   ,16'd8856};
dout[132]={ 4'd5     ,  4'd6, 16'd54908   ,16'd10627};
dout[133]={ 4'd5     ,  4'd6, 16'd53137   ,16'd12398};
dout[134]={ 4'd5     ,  4'd6, 16'd51366   ,16'd14169};
dout[135]={ 4'd5     ,  4'd6, 16'd49594   ,16'd15941};
dout[136]={ 4'd5     ,  4'd6, 16'd47823   ,16'd17712};
dout[137]={ 4'd5     ,  4'd6, 16'd46052   ,16'd19483};
dout[138]={ 4'd5     ,  4'd6, 16'd44281   ,16'd21254};
dout[139]={ 4'd5     ,  4'd6, 16'd42509   ,16'd23026};
dout[140]={ 4'd5     ,  4'd6, 16'd40738   ,16'd24797};
dout[141]={ 4'd5     ,  4'd6, 16'd38967   ,16'd26568};
dout[142]={ 4'd5     ,  4'd6, 16'd37196   ,16'd28339};
dout[143]={ 4'd5     ,  4'd6, 16'd35424   ,16'd30111};
dout[144]={ 4'd5     ,  4'd6, 16'd33653   ,16'd31882};
dout[145]={ 4'd5     ,  4'd6, 16'd31882   ,16'd33653};
dout[146]={ 4'd5     ,  4'd6, 16'd30111   ,16'd35424};
dout[147]={ 4'd5     ,  4'd6, 16'd28339   ,16'd37196};
dout[148]={ 4'd5     ,  4'd6, 16'd26568   ,16'd38967};
dout[149]={ 4'd5     ,  4'd6, 16'd24797   ,16'd40738};
dout[150]={ 4'd5     ,  4'd6, 16'd23026   ,16'd42509};
dout[151]={ 4'd5     ,  4'd6, 16'd21254   ,16'd44281};
dout[152]={ 4'd5     ,  4'd6, 16'd19483   ,16'd46052};
dout[153]={ 4'd5     ,  4'd6, 16'd17712   ,16'd47823};
dout[154]={ 4'd5     ,  4'd6, 16'd15941   ,16'd49594};
dout[155]={ 4'd5     ,  4'd6, 16'd14169   ,16'd51366};
dout[156]={ 4'd5     ,  4'd6, 16'd12398   ,16'd53137};
dout[157]={ 4'd5     ,  4'd6, 16'd10627   ,16'd54908};
dout[158]={ 4'd5     ,  4'd6, 16'd8856   ,16'd56679};
dout[159]={ 4'd5     ,  4'd6, 16'd7084   ,16'd58451};
dout[160]={ 4'd5     ,  4'd6, 16'd5313   ,16'd60222};
dout[161]={ 4'd5     ,  4'd6, 16'd3542   ,16'd61993};
dout[162]={ 4'd5     ,  4'd6, 16'd1771   ,16'd63764};
dout[163]={ 4'd6     ,  4'd0, 16'd65535   ,16'd0};
dout[164]={ 4'd6     ,  4'd7, 16'd64079   ,16'd1456};
dout[165]={ 4'd6     ,  4'd7, 16'd62623   ,16'd2912};
dout[166]={ 4'd6     ,  4'd7, 16'd61166   ,16'd4369};
dout[167]={ 4'd6     ,  4'd7, 16'd59710   ,16'd5825};
dout[168]={ 4'd6     ,  4'd7, 16'd58254   ,16'd7281};
dout[169]={ 4'd6     ,  4'd7, 16'd56797   ,16'd8738};
dout[170]={ 4'd6     ,  4'd7, 16'd55341   ,16'd10194};
dout[171]={ 4'd6     ,  4'd7, 16'd53885   ,16'd11650};
dout[172]={ 4'd6     ,  4'd7, 16'd52428   ,16'd13107};
dout[173]={ 4'd6     ,  4'd7, 16'd50972   ,16'd14563};
dout[174]={ 4'd6     ,  4'd7, 16'd49516   ,16'd16019};
dout[175]={ 4'd6     ,  4'd7, 16'd48059   ,16'd17476};
dout[176]={ 4'd6     ,  4'd7, 16'd46603   ,16'd18932};
dout[177]={ 4'd6     ,  4'd7, 16'd45147   ,16'd20388};
dout[178]={ 4'd6     ,  4'd7, 16'd43690   ,16'd21845};
dout[179]={ 4'd6     ,  4'd7, 16'd42234   ,16'd23301};
dout[180]={ 4'd6     ,  4'd7, 16'd40777   ,16'd24758};
dout[181]={ 4'd6     ,  4'd7, 16'd39321   ,16'd26214};
dout[182]={ 4'd6     ,  4'd7, 16'd37865   ,16'd27670};
dout[183]={ 4'd6     ,  4'd7, 16'd36408   ,16'd29127};
dout[184]={ 4'd6     ,  4'd7, 16'd34952   ,16'd30583};
dout[185]={ 4'd6     ,  4'd7, 16'd33496   ,16'd32039};
dout[186]={ 4'd6     ,  4'd7, 16'd32039   ,16'd33496};
dout[187]={ 4'd6     ,  4'd7, 16'd30583   ,16'd34952};
dout[188]={ 4'd6     ,  4'd7, 16'd29127   ,16'd36408};
dout[189]={ 4'd6     ,  4'd7, 16'd27670   ,16'd37865};
dout[190]={ 4'd6     ,  4'd7, 16'd26214   ,16'd39321};
dout[191]={ 4'd6     ,  4'd7, 16'd24758   ,16'd40777};
dout[192]={ 4'd6     ,  4'd7, 16'd23301   ,16'd42234};
dout[193]={ 4'd6     ,  4'd7, 16'd21845   ,16'd43690};
dout[194]={ 4'd6     ,  4'd7, 16'd20388   ,16'd45147};
dout[195]={ 4'd6     ,  4'd7, 16'd18932   ,16'd46603};
dout[196]={ 4'd6     ,  4'd7, 16'd17476   ,16'd48059};
dout[197]={ 4'd6     ,  4'd7, 16'd16019   ,16'd49516};
dout[198]={ 4'd6     ,  4'd7, 16'd14563   ,16'd50972};
dout[199]={ 4'd6     ,  4'd7, 16'd13107   ,16'd52428};
dout[200]={ 4'd6     ,  4'd7, 16'd11650   ,16'd53885};
dout[201]={ 4'd6     ,  4'd7, 16'd10194   ,16'd55341};
dout[202]={ 4'd6     ,  4'd7, 16'd8738   ,16'd56797};
dout[203]={ 4'd6     ,  4'd7, 16'd7281   ,16'd58254};
dout[204]={ 4'd6     ,  4'd7, 16'd5825   ,16'd59710};
dout[205]={ 4'd6     ,  4'd7, 16'd4369   ,16'd61166};
dout[206]={ 4'd6     ,  4'd7, 16'd2912   ,16'd62623};
dout[207]={ 4'd6     ,  4'd7, 16'd1456   ,16'd64079};
dout[208]={ 4'd7     ,  4'd0, 16'd65535   ,16'd0};
dout[209]={ 4'd7     ,  4'd8, 16'd64365   ,16'd1170};
dout[210]={ 4'd7     ,  4'd8, 16'd63195   ,16'd2340};
dout[211]={ 4'd7     ,  4'd8, 16'd62025   ,16'd3510};
dout[212]={ 4'd7     ,  4'd8, 16'd60854   ,16'd4681};
dout[213]={ 4'd7     ,  4'd8, 16'd59684   ,16'd5851};
dout[214]={ 4'd7     ,  4'd8, 16'd58514   ,16'd7021};
dout[215]={ 4'd7     ,  4'd8, 16'd57344   ,16'd8192};
dout[216]={ 4'd7     ,  4'd8, 16'd56173   ,16'd9362};
dout[217]={ 4'd7     ,  4'd8, 16'd55003   ,16'd10532};
dout[218]={ 4'd7     ,  4'd8, 16'd53833   ,16'd11702};
dout[219]={ 4'd7     ,  4'd8, 16'd52662   ,16'd12873};
dout[220]={ 4'd7     ,  4'd8, 16'd51492   ,16'd14043};
dout[221]={ 4'd7     ,  4'd8, 16'd50322   ,16'd15213};
dout[222]={ 4'd7     ,  4'd8, 16'd49152   ,16'd16384};
dout[223]={ 4'd7     ,  4'd8, 16'd47981   ,16'd17554};
dout[224]={ 4'd7     ,  4'd8, 16'd46811   ,16'd18724};
dout[225]={ 4'd7     ,  4'd8, 16'd45641   ,16'd19894};
dout[226]={ 4'd7     ,  4'd8, 16'd44470   ,16'd21065};
dout[227]={ 4'd7     ,  4'd8, 16'd43300   ,16'd22235};
dout[228]={ 4'd7     ,  4'd8, 16'd42130   ,16'd23405};
dout[229]={ 4'd7     ,  4'd8, 16'd40960   ,16'd24576};
dout[230]={ 4'd7     ,  4'd8, 16'd39789   ,16'd25746};
dout[231]={ 4'd7     ,  4'd8, 16'd38619   ,16'd26916};
dout[232]={ 4'd7     ,  4'd8, 16'd37449   ,16'd28086};
dout[233]={ 4'd7     ,  4'd8, 16'd36278   ,16'd29257};
dout[234]={ 4'd7     ,  4'd8, 16'd35108   ,16'd30427};
dout[235]={ 4'd7     ,  4'd8, 16'd33938   ,16'd31597};
dout[236]={ 4'd7     ,  4'd8, 16'd32768   ,16'd32768};
dout[237]={ 4'd7     ,  4'd8, 16'd31597   ,16'd33938};
dout[238]={ 4'd7     ,  4'd8, 16'd30427   ,16'd35108};
dout[239]={ 4'd7     ,  4'd8, 16'd29257   ,16'd36278};
dout[240]={ 4'd7     ,  4'd8, 16'd28086   ,16'd37449};
dout[241]={ 4'd7     ,  4'd8, 16'd26916   ,16'd38619};
dout[242]={ 4'd7     ,  4'd8, 16'd25746   ,16'd39789};
dout[243]={ 4'd7     ,  4'd8, 16'd24576   ,16'd40960};
dout[244]={ 4'd7     ,  4'd8, 16'd23405   ,16'd42130};
dout[245]={ 4'd7     ,  4'd8, 16'd22235   ,16'd43300};
dout[246]={ 4'd7     ,  4'd8, 16'd21065   ,16'd44470};
dout[247]={ 4'd7     ,  4'd8, 16'd19894   ,16'd45641};
dout[248]={ 4'd7     ,  4'd8, 16'd18724   ,16'd46811};
dout[249]={ 4'd7     ,  4'd8, 16'd17554   ,16'd47981};
dout[250]={ 4'd7     ,  4'd8, 16'd16384   ,16'd49152};
dout[251]={ 4'd7     ,  4'd8, 16'd15213   ,16'd50322};
dout[252]={ 4'd7     ,  4'd8, 16'd14043   ,16'd51492};
dout[253]={ 4'd7     ,  4'd8, 16'd12873   ,16'd52662};
dout[254]={ 4'd7     ,  4'd8, 16'd11702   ,16'd53833};
dout[255]={ 4'd7     ,  4'd8, 16'd10532   ,16'd55003};
dout[256]={ 4'd7     ,  4'd8, 16'd9362   ,16'd56173};
dout[257]={ 4'd7     ,  4'd8, 16'd8192   ,16'd57344};
dout[258]={ 4'd7     ,  4'd8, 16'd7021   ,16'd58514};
dout[259]={ 4'd7     ,  4'd8, 16'd5851   ,16'd59684};
dout[260]={ 4'd7     ,  4'd8, 16'd4681   ,16'd60854};
dout[261]={ 4'd7     ,  4'd8, 16'd3510   ,16'd62025};
dout[262]={ 4'd7     ,  4'd8, 16'd2340   ,16'd63195};
dout[263]={ 4'd7     ,  4'd8, 16'd1170   ,16'd64365};
dout[264]={ 4'd8     ,  4'd0, 16'd65535   ,16'd0};
dout[265]={ 4'd8     ,  4'd9, 16'd64557   ,16'd978};
dout[266]={ 4'd8     ,  4'd9, 16'd63579   ,16'd1956};
dout[267]={ 4'd8     ,  4'd9, 16'd62601   ,16'd2934};
dout[268]={ 4'd8     ,  4'd9, 16'd61623   ,16'd3912};
dout[269]={ 4'd8     ,  4'd9, 16'd60645   ,16'd4890};
dout[270]={ 4'd8     ,  4'd9, 16'd59667   ,16'd5868};
dout[271]={ 4'd8     ,  4'd9, 16'd58688   ,16'd6847};
dout[272]={ 4'd8     ,  4'd9, 16'd57710   ,16'd7825};
dout[273]={ 4'd8     ,  4'd9, 16'd56732   ,16'd8803};
dout[274]={ 4'd8     ,  4'd9, 16'd55754   ,16'd9781};
dout[275]={ 4'd8     ,  4'd9, 16'd54776   ,16'd10759};
dout[276]={ 4'd8     ,  4'd9, 16'd53798   ,16'd11737};
dout[277]={ 4'd8     ,  4'd9, 16'd52820   ,16'd12715};
dout[278]={ 4'd8     ,  4'd9, 16'd51841   ,16'd13694};
dout[279]={ 4'd8     ,  4'd9, 16'd50863   ,16'd14672};
dout[280]={ 4'd8     ,  4'd9, 16'd49885   ,16'd15650};
dout[281]={ 4'd8     ,  4'd9, 16'd48907   ,16'd16628};
dout[282]={ 4'd8     ,  4'd9, 16'd47929   ,16'd17606};
dout[283]={ 4'd8     ,  4'd9, 16'd46951   ,16'd18584};
dout[284]={ 4'd8     ,  4'd9, 16'd45973   ,16'd19562};
dout[285]={ 4'd8     ,  4'd9, 16'd44994   ,16'd20541};
dout[286]={ 4'd8     ,  4'd9, 16'd44016   ,16'd21519};
dout[287]={ 4'd8     ,  4'd9, 16'd43038   ,16'd22497};
dout[288]={ 4'd8     ,  4'd9, 16'd42060   ,16'd23475};
dout[289]={ 4'd8     ,  4'd9, 16'd41082   ,16'd24453};
dout[290]={ 4'd8     ,  4'd9, 16'd40104   ,16'd25431};
dout[291]={ 4'd8     ,  4'd9, 16'd39125   ,16'd26410};
dout[292]={ 4'd8     ,  4'd9, 16'd38147   ,16'd27388};
dout[293]={ 4'd8     ,  4'd9, 16'd37169   ,16'd28366};
dout[294]={ 4'd8     ,  4'd9, 16'd36191   ,16'd29344};
dout[295]={ 4'd8     ,  4'd9, 16'd35213   ,16'd30322};
dout[296]={ 4'd8     ,  4'd9, 16'd34235   ,16'd31300};
dout[297]={ 4'd8     ,  4'd9, 16'd33257   ,16'd32278};
dout[298]={ 4'd8     ,  4'd9, 16'd32278   ,16'd33257};
dout[299]={ 4'd8     ,  4'd9, 16'd31300   ,16'd34235};
dout[300]={ 4'd8     ,  4'd9, 16'd30322   ,16'd35213};
dout[301]={ 4'd8     ,  4'd9, 16'd29344   ,16'd36191};
dout[302]={ 4'd8     ,  4'd9, 16'd28366   ,16'd37169};
dout[303]={ 4'd8     ,  4'd9, 16'd27388   ,16'd38147};
dout[304]={ 4'd8     ,  4'd9, 16'd26410   ,16'd39125};
dout[305]={ 4'd8     ,  4'd9, 16'd25431   ,16'd40104};
dout[306]={ 4'd8     ,  4'd9, 16'd24453   ,16'd41082};
dout[307]={ 4'd8     ,  4'd9, 16'd23475   ,16'd42060};
dout[308]={ 4'd8     ,  4'd9, 16'd22497   ,16'd43038};
dout[309]={ 4'd8     ,  4'd9, 16'd21519   ,16'd44016};
dout[310]={ 4'd8     ,  4'd9, 16'd20541   ,16'd44994};
dout[311]={ 4'd8     ,  4'd9, 16'd19562   ,16'd45973};
dout[312]={ 4'd8     ,  4'd9, 16'd18584   ,16'd46951};
dout[313]={ 4'd8     ,  4'd9, 16'd17606   ,16'd47929};
dout[314]={ 4'd8     ,  4'd9, 16'd16628   ,16'd48907};
dout[315]={ 4'd8     ,  4'd9, 16'd15650   ,16'd49885};
dout[316]={ 4'd8     ,  4'd9, 16'd14672   ,16'd50863};
dout[317]={ 4'd8     ,  4'd9, 16'd13694   ,16'd51841};
dout[318]={ 4'd8     ,  4'd9, 16'd12715   ,16'd52820};
dout[319]={ 4'd8     ,  4'd9, 16'd11737   ,16'd53798};
dout[320]={ 4'd8     ,  4'd9, 16'd10759   ,16'd54776};
dout[321]={ 4'd8     ,  4'd9, 16'd9781   ,16'd55754};
dout[322]={ 4'd8     ,  4'd9, 16'd8803   ,16'd56732};
dout[323]={ 4'd8     ,  4'd9, 16'd7825   ,16'd57710};
dout[324]={ 4'd8     ,  4'd9, 16'd6847   ,16'd58688};
dout[325]={ 4'd8     ,  4'd9, 16'd5868   ,16'd59667};
dout[326]={ 4'd8     ,  4'd9, 16'd4890   ,16'd60645};
dout[327]={ 4'd8     ,  4'd9, 16'd3912   ,16'd61623};
dout[328]={ 4'd8     ,  4'd9, 16'd2934   ,16'd62601};
dout[329]={ 4'd8     ,  4'd9, 16'd1956   ,16'd63579};
dout[330]={ 4'd8     ,  4'd9, 16'd978   ,16'd64557};
dout[331]={ 4'd9     ,  4'd0, 16'd65535   ,16'd0};
dout[332]={ 4'd9     ,  4'd10, 16'd64726   ,16'd809};
dout[333]={ 4'd9     ,  4'd10, 16'd63917   ,16'd1618};
dout[334]={ 4'd9     ,  4'd10, 16'd63108   ,16'd2427};
dout[335]={ 4'd9     ,  4'd10, 16'd62299   ,16'd3236};
dout[336]={ 4'd9     ,  4'd10, 16'd61490   ,16'd4045};
dout[337]={ 4'd9     ,  4'd10, 16'd60681   ,16'd4854};
dout[338]={ 4'd9     ,  4'd10, 16'd59872   ,16'd5663};
dout[339]={ 4'd9     ,  4'd10, 16'd59063   ,16'd6472};
dout[340]={ 4'd9     ,  4'd10, 16'd58254   ,16'd7281};
dout[341]={ 4'd9     ,  4'd10, 16'd57445   ,16'd8090};
dout[342]={ 4'd9     ,  4'd10, 16'd56636   ,16'd8899};
dout[343]={ 4'd9     ,  4'd10, 16'd55826   ,16'd9709};
dout[344]={ 4'd9     ,  4'd10, 16'd55017   ,16'd10518};
dout[345]={ 4'd9     ,  4'd10, 16'd54208   ,16'd11327};
dout[346]={ 4'd9     ,  4'd10, 16'd53399   ,16'd12136};
dout[347]={ 4'd9     ,  4'd10, 16'd52590   ,16'd12945};
dout[348]={ 4'd9     ,  4'd10, 16'd51781   ,16'd13754};
dout[349]={ 4'd9     ,  4'd10, 16'd50972   ,16'd14563};
dout[350]={ 4'd9     ,  4'd10, 16'd50163   ,16'd15372};
dout[351]={ 4'd9     ,  4'd10, 16'd49354   ,16'd16181};
dout[352]={ 4'd9     ,  4'd10, 16'd48545   ,16'd16990};
dout[353]={ 4'd9     ,  4'd10, 16'd47736   ,16'd17799};
dout[354]={ 4'd9     ,  4'd10, 16'd46927   ,16'd18608};
dout[355]={ 4'd9     ,  4'd10, 16'd46117   ,16'd19418};
dout[356]={ 4'd9     ,  4'd10, 16'd45308   ,16'd20227};
dout[357]={ 4'd9     ,  4'd10, 16'd44499   ,16'd21036};
dout[358]={ 4'd9     ,  4'd10, 16'd43690   ,16'd21845};
dout[359]={ 4'd9     ,  4'd10, 16'd42881   ,16'd22654};
dout[360]={ 4'd9     ,  4'd10, 16'd42072   ,16'd23463};
dout[361]={ 4'd9     ,  4'd10, 16'd41263   ,16'd24272};
dout[362]={ 4'd9     ,  4'd10, 16'd40454   ,16'd25081};
dout[363]={ 4'd9     ,  4'd10, 16'd39645   ,16'd25890};
dout[364]={ 4'd9     ,  4'd10, 16'd38836   ,16'd26699};
dout[365]={ 4'd9     ,  4'd10, 16'd38027   ,16'd27508};
dout[366]={ 4'd9     ,  4'd10, 16'd37217   ,16'd28318};
dout[367]={ 4'd9     ,  4'd10, 16'd36408   ,16'd29127};
dout[368]={ 4'd9     ,  4'd10, 16'd35599   ,16'd29936};
dout[369]={ 4'd9     ,  4'd10, 16'd34790   ,16'd30745};
dout[370]={ 4'd9     ,  4'd10, 16'd33981   ,16'd31554};
dout[371]={ 4'd9     ,  4'd10, 16'd33172   ,16'd32363};
dout[372]={ 4'd9     ,  4'd10, 16'd32363   ,16'd33172};
dout[373]={ 4'd9     ,  4'd10, 16'd31554   ,16'd33981};
dout[374]={ 4'd9     ,  4'd10, 16'd30745   ,16'd34790};
dout[375]={ 4'd9     ,  4'd10, 16'd29936   ,16'd35599};
dout[376]={ 4'd9     ,  4'd10, 16'd29127   ,16'd36408};
dout[377]={ 4'd9     ,  4'd10, 16'd28318   ,16'd37217};
dout[378]={ 4'd9     ,  4'd10, 16'd27508   ,16'd38027};
dout[379]={ 4'd9     ,  4'd10, 16'd26699   ,16'd38836};
dout[380]={ 4'd9     ,  4'd10, 16'd25890   ,16'd39645};
dout[381]={ 4'd9     ,  4'd10, 16'd25081   ,16'd40454};
dout[382]={ 4'd9     ,  4'd10, 16'd24272   ,16'd41263};
dout[383]={ 4'd9     ,  4'd10, 16'd23463   ,16'd42072};
dout[384]={ 4'd9     ,  4'd10, 16'd22654   ,16'd42881};
dout[385]={ 4'd9     ,  4'd10, 16'd21845   ,16'd43690};
dout[386]={ 4'd9     ,  4'd10, 16'd21036   ,16'd44499};
dout[387]={ 4'd9     ,  4'd10, 16'd20227   ,16'd45308};
dout[388]={ 4'd9     ,  4'd10, 16'd19418   ,16'd46117};
dout[389]={ 4'd9     ,  4'd10, 16'd18608   ,16'd46927};
dout[390]={ 4'd9     ,  4'd10, 16'd17799   ,16'd47736};
dout[391]={ 4'd9     ,  4'd10, 16'd16990   ,16'd48545};
dout[392]={ 4'd9     ,  4'd10, 16'd16181   ,16'd49354};
dout[393]={ 4'd9     ,  4'd10, 16'd15372   ,16'd50163};
dout[394]={ 4'd9     ,  4'd10, 16'd14563   ,16'd50972};
dout[395]={ 4'd9     ,  4'd10, 16'd13754   ,16'd51781};
dout[396]={ 4'd9     ,  4'd10, 16'd12945   ,16'd52590};
dout[397]={ 4'd9     ,  4'd10, 16'd12136   ,16'd53399};
dout[398]={ 4'd9     ,  4'd10, 16'd11327   ,16'd54208};
dout[399]={ 4'd9     ,  4'd10, 16'd10518   ,16'd55017};
dout[400]={ 4'd9     ,  4'd10, 16'd9709   ,16'd55826};
dout[401]={ 4'd9     ,  4'd10, 16'd8899   ,16'd56636};
dout[402]={ 4'd9     ,  4'd10, 16'd8090   ,16'd57445};
dout[403]={ 4'd9     ,  4'd10, 16'd7281   ,16'd58254};
dout[404]={ 4'd9     ,  4'd10, 16'd6472   ,16'd59063};
dout[405]={ 4'd9     ,  4'd10, 16'd5663   ,16'd59872};
dout[406]={ 4'd9     ,  4'd10, 16'd4854   ,16'd60681};
dout[407]={ 4'd9     ,  4'd10, 16'd4045   ,16'd61490};
dout[408]={ 4'd9     ,  4'd10, 16'd3236   ,16'd62299};
dout[409]={ 4'd9     ,  4'd10, 16'd2427   ,16'd63108};
dout[410]={ 4'd9     ,  4'd10, 16'd1618   ,16'd63917};
dout[411]={ 4'd9     ,  4'd10, 16'd809   ,16'd64726};
dout[412]={ 4'd10     ,  4'd0, 16'd65535   ,16'd0};
dout[413]={ 4'd10     ,  4'd0, 16'd64880   ,16'd0};
dout[414]={ 4'd10     ,  4'd0, 16'd64225   ,16'd0};
dout[415]={ 4'd10     ,  4'd0, 16'd63569   ,16'd0};
dout[416]={ 4'd10     ,  4'd0, 16'd62914   ,16'd0};
dout[417]={ 4'd10     ,  4'd0, 16'd62259   ,16'd0};
dout[418]={ 4'd10     ,  4'd0, 16'd61603   ,16'd0};
dout[419]={ 4'd10     ,  4'd0, 16'd60948   ,16'd0};
dout[420]={ 4'd10     ,  4'd0, 16'd60293   ,16'd0};
dout[421]={ 4'd10     ,  4'd0, 16'd59637   ,16'd0};
dout[422]={ 4'd10     ,  4'd0, 16'd58982   ,16'd0};
dout[423]={ 4'd10     ,  4'd0, 16'd58327   ,16'd0};
dout[424]={ 4'd10     ,  4'd0, 16'd57671   ,16'd0};
dout[425]={ 4'd10     ,  4'd0, 16'd57016   ,16'd0};
dout[426]={ 4'd10     ,  4'd0, 16'd56360   ,16'd0};
dout[427]={ 4'd10     ,  4'd0, 16'd55705   ,16'd0};
dout[428]={ 4'd10     ,  4'd0, 16'd55050   ,16'd0};
dout[429]={ 4'd10     ,  4'd0, 16'd54394   ,16'd0};
dout[430]={ 4'd10     ,  4'd0, 16'd53739   ,16'd0};
dout[431]={ 4'd10     ,  4'd0, 16'd53084   ,16'd0};
dout[432]={ 4'd10     ,  4'd0, 16'd52428   ,16'd0};
dout[433]={ 4'd10     ,  4'd0, 16'd51773   ,16'd0};
dout[434]={ 4'd10     ,  4'd0, 16'd51118   ,16'd0};
dout[435]={ 4'd10     ,  4'd0, 16'd50462   ,16'd0};
dout[436]={ 4'd10     ,  4'd0, 16'd49807   ,16'd0};
dout[437]={ 4'd10     ,  4'd0, 16'd49152   ,16'd0};
dout[438]={ 4'd10     ,  4'd0, 16'd48496   ,16'd0};
dout[439]={ 4'd10     ,  4'd0, 16'd47841   ,16'd0};
dout[440]={ 4'd10     ,  4'd0, 16'd47185   ,16'd0};
dout[441]={ 4'd10     ,  4'd0, 16'd46530   ,16'd0};
dout[442]={ 4'd10     ,  4'd0, 16'd45875   ,16'd0};
dout[443]={ 4'd10     ,  4'd0, 16'd45219   ,16'd0};
dout[444]={ 4'd10     ,  4'd0, 16'd44564   ,16'd0};
dout[445]={ 4'd10     ,  4'd0, 16'd43909   ,16'd0};
dout[446]={ 4'd10     ,  4'd0, 16'd43253   ,16'd0};
dout[447]={ 4'd10     ,  4'd0, 16'd42598   ,16'd0};
dout[448]={ 4'd10     ,  4'd0, 16'd41943   ,16'd0};
dout[449]={ 4'd10     ,  4'd0, 16'd41287   ,16'd0};
dout[450]={ 4'd10     ,  4'd0, 16'd40632   ,16'd0};
dout[451]={ 4'd10     ,  4'd0, 16'd39976   ,16'd0};
dout[452]={ 4'd10     ,  4'd0, 16'd39321   ,16'd0};
dout[453]={ 4'd10     ,  4'd0, 16'd38666   ,16'd0};
dout[454]={ 4'd10     ,  4'd0, 16'd38010   ,16'd0};
dout[455]={ 4'd10     ,  4'd0, 16'd37355   ,16'd0};
dout[456]={ 4'd10     ,  4'd0, 16'd36700   ,16'd0};
dout[457]={ 4'd10     ,  4'd0, 16'd36044   ,16'd0};
dout[458]={ 4'd10     ,  4'd0, 16'd35389   ,16'd0};
dout[459]={ 4'd10     ,  4'd0, 16'd34734   ,16'd0};
dout[460]={ 4'd10     ,  4'd0, 16'd34078   ,16'd0};
dout[461]={ 4'd10     ,  4'd0, 16'd33423   ,16'd0};
dout[462]={ 4'd10     ,  4'd0, 16'd32768   ,16'd0};
dout[463]={ 4'd10     ,  4'd0, 16'd32112   ,16'd0};
dout[464]={ 4'd10     ,  4'd0, 16'd31457   ,16'd0};
dout[465]={ 4'd10     ,  4'd0, 16'd30801   ,16'd0};
dout[466]={ 4'd10     ,  4'd0, 16'd30146   ,16'd0};
dout[467]={ 4'd10     ,  4'd0, 16'd29491   ,16'd0};
dout[468]={ 4'd10     ,  4'd0, 16'd28835   ,16'd0};
dout[469]={ 4'd10     ,  4'd0, 16'd28180   ,16'd0};
dout[470]={ 4'd10     ,  4'd0, 16'd27525   ,16'd0};
dout[471]={ 4'd10     ,  4'd0, 16'd26869   ,16'd0};
dout[472]={ 4'd10     ,  4'd0, 16'd26214   ,16'd0};
dout[473]={ 4'd10     ,  4'd0, 16'd25559   ,16'd0};
dout[474]={ 4'd10     ,  4'd0, 16'd24903   ,16'd0};
dout[475]={ 4'd10     ,  4'd0, 16'd24248   ,16'd0};
dout[476]={ 4'd10     ,  4'd0, 16'd23592   ,16'd0};
dout[477]={ 4'd10     ,  4'd0, 16'd22937   ,16'd0};
dout[478]={ 4'd10     ,  4'd0, 16'd22282   ,16'd0};
dout[479]={ 4'd10     ,  4'd0, 16'd21626   ,16'd0};
dout[480]={ 4'd10     ,  4'd0, 16'd20971   ,16'd0};
dout[481]={ 4'd10     ,  4'd0, 16'd20316   ,16'd0};
dout[482]={ 4'd10     ,  4'd0, 16'd19660   ,16'd0};
dout[483]={ 4'd10     ,  4'd0, 16'd19005   ,16'd0};
dout[484]={ 4'd10     ,  4'd0, 16'd18350   ,16'd0};
dout[485]={ 4'd10     ,  4'd0, 16'd17694   ,16'd0};
dout[486]={ 4'd10     ,  4'd0, 16'd17039   ,16'd0};
dout[487]={ 4'd10     ,  4'd0, 16'd16384   ,16'd0};
dout[488]={ 4'd10     ,  4'd0, 16'd15728   ,16'd0};
dout[489]={ 4'd10     ,  4'd0, 16'd15073   ,16'd0};
dout[490]={ 4'd10     ,  4'd0, 16'd14417   ,16'd0};
dout[491]={ 4'd10     ,  4'd0, 16'd13762   ,16'd0};
dout[492]={ 4'd10     ,  4'd0, 16'd13107   ,16'd0};
dout[493]={ 4'd10     ,  4'd0, 16'd12451   ,16'd0};
dout[494]={ 4'd10     ,  4'd0, 16'd11796   ,16'd0};
dout[495]={ 4'd10     ,  4'd0, 16'd11141   ,16'd0};
dout[496]={ 4'd10     ,  4'd0, 16'd10485   ,16'd0};
dout[497]={ 4'd10     ,  4'd0, 16'd9830   ,16'd0};
dout[498]={ 4'd10     ,  4'd0, 16'd9175   ,16'd0};
dout[499]={ 4'd10     ,  4'd0, 16'd8519   ,16'd0};
dout[500]={ 4'd10     ,  4'd0, 16'd7864   ,16'd0};
dout[501]={ 4'd10     ,  4'd0, 16'd7208   ,16'd0};
dout[502]={ 4'd10     ,  4'd0, 16'd6553   ,16'd0};
dout[503]={ 4'd10     ,  4'd0, 16'd5898   ,16'd0};
dout[504]={ 4'd10     ,  4'd0, 16'd5242   ,16'd0};
dout[505]={ 4'd10     ,  4'd0, 16'd4587   ,16'd0};
dout[506]={ 4'd10     ,  4'd0, 16'd3932   ,16'd0};
dout[507]={ 4'd10     ,  4'd0, 16'd3276   ,16'd0};
dout[508]={ 4'd10     ,  4'd0, 16'd2621   ,16'd0};
dout[509]={ 4'd10     ,  4'd0, 16'd1966   ,16'd0};
dout[510]={ 4'd10     ,  4'd0, 16'd1310   ,16'd0};
dout[511]={ 4'd10     ,  4'd0, 16'd655   ,16'd0};
dout[512]={ 4'd0     ,  4'd0, 16'd0   ,16'd0};
dout[513]=40'b0;
dout[514]=40'b0;
dout[515]=40'b0;
dout[516]=40'b0;
dout[517]=40'b0;
dout[518]=40'b0;
dout[519]=40'b0;
dout[520]=40'b0;
dout[521]=40'b0;
dout[522]=40'b0;
dout[523]=40'b0;
dout[524]=40'b0;
dout[525]=40'b0;
dout[526]=40'b0;
dout[527]=40'b0;
dout[528]=40'b0;
dout[529]=40'b0;
dout[530]=40'b0;
dout[531]=40'b0;
dout[532]=40'b0;
dout[533]=40'b0;
dout[534]=40'b0;
dout[535]=40'b0;
dout[536]=40'b0;
dout[537]=40'b0;
dout[538]=40'b0;
dout[539]=40'b0;
dout[540]=40'b0;
dout[541]=40'b0;
dout[542]=40'b0;
dout[543]=40'b0;
dout[544]=40'b0;
dout[545]=40'b0;
dout[546]=40'b0;
dout[547]=40'b0;
dout[548]=40'b0;
dout[549]=40'b0;
dout[550]=40'b0;
dout[551]=40'b0;
dout[552]=40'b0;
dout[553]=40'b0;
dout[554]=40'b0;
dout[555]=40'b0;
dout[556]=40'b0;
dout[557]=40'b0;
dout[558]=40'b0;
dout[559]=40'b0;
dout[560]=40'b0;
dout[561]=40'b0;
dout[562]=40'b0;
dout[563]=40'b0;
dout[564]=40'b0;
dout[565]=40'b0;
dout[566]=40'b0;
dout[567]=40'b0;
dout[568]=40'b0;
dout[569]=40'b0;
dout[570]=40'b0;
dout[571]=40'b0;
dout[572]=40'b0;
dout[573]=40'b0;
dout[574]=40'b0;
dout[575]=40'b0;
dout[576]=40'b0;
dout[577]=40'b0;
dout[578]=40'b0;
dout[579]=40'b0;
dout[580]=40'b0;
dout[581]=40'b0;
dout[582]=40'b0;
dout[583]=40'b0;
dout[584]=40'b0;
dout[585]=40'b0;
dout[586]=40'b0;
dout[587]=40'b0;
dout[588]=40'b0;
dout[589]=40'b0;
dout[590]=40'b0;
dout[591]=40'b0;
dout[592]=40'b0;
dout[593]=40'b0;
dout[594]=40'b0;
dout[595]=40'b0;
dout[596]=40'b0;
dout[597]=40'b0;
dout[598]=40'b0;
dout[599]=40'b0;
dout[600]=40'b0;
dout[601]=40'b0;
dout[602]=40'b0;
dout[603]=40'b0;
dout[604]=40'b0;
dout[605]=40'b0;
dout[606]=40'b0;
dout[607]=40'b0;
dout[608]=40'b0;
dout[609]=40'b0;
dout[610]=40'b0;
dout[611]=40'b0;
dout[612]=40'b0;
dout[613]=40'b0;
dout[614]=40'b0;
dout[615]=40'b0;
dout[616]=40'b0;
dout[617]=40'b0;
dout[618]=40'b0;
dout[619]=40'b0;
dout[620]=40'b0;
dout[621]=40'b0;
dout[622]=40'b0;
dout[623]=40'b0;
dout[624]=40'b0;
dout[625]=40'b0;
dout[626]=40'b0;
dout[627]=40'b0;
dout[628]=40'b0;
dout[629]=40'b0;
dout[630]=40'b0;
dout[631]=40'b0;
dout[632]=40'b0;
dout[633]=40'b0;
dout[634]=40'b0;
dout[635]=40'b0;
dout[636]=40'b0;
dout[637]=40'b0;
dout[638]=40'b0;
dout[639]=40'b0;
dout[640]=40'b0;
dout[641]=40'b0;
dout[642]=40'b0;
dout[643]=40'b0;
dout[644]=40'b0;
dout[645]=40'b0;
dout[646]=40'b0;
dout[647]=40'b0;
dout[648]=40'b0;
dout[649]=40'b0;
dout[650]=40'b0;
dout[651]=40'b0;
dout[652]=40'b0;
dout[653]=40'b0;
dout[654]=40'b0;
dout[655]=40'b0;
dout[656]=40'b0;
dout[657]=40'b0;
dout[658]=40'b0;
dout[659]=40'b0;
dout[660]=40'b0;
dout[661]=40'b0;
dout[662]=40'b0;
dout[663]=40'b0;
dout[664]=40'b0;
dout[665]=40'b0;
dout[666]=40'b0;
dout[667]=40'b0;
dout[668]=40'b0;
dout[669]=40'b0;
dout[670]=40'b0;
dout[671]=40'b0;
dout[672]=40'b0;
dout[673]=40'b0;
dout[674]=40'b0;
dout[675]=40'b0;
dout[676]=40'b0;
dout[677]=40'b0;
dout[678]=40'b0;
dout[679]=40'b0;
dout[680]=40'b0;
dout[681]=40'b0;
dout[682]=40'b0;
dout[683]=40'b0;
dout[684]=40'b0;
dout[685]=40'b0;
dout[686]=40'b0;
dout[687]=40'b0;
dout[688]=40'b0;
dout[689]=40'b0;
dout[690]=40'b0;
dout[691]=40'b0;
dout[692]=40'b0;
dout[693]=40'b0;
dout[694]=40'b0;
dout[695]=40'b0;
dout[696]=40'b0;
dout[697]=40'b0;
dout[698]=40'b0;
dout[699]=40'b0;
dout[700]=40'b0;
dout[701]=40'b0;
dout[702]=40'b0;
dout[703]=40'b0;
dout[704]=40'b0;
dout[705]=40'b0;
dout[706]=40'b0;
dout[707]=40'b0;
dout[708]=40'b0;
dout[709]=40'b0;
dout[710]=40'b0;
dout[711]=40'b0;
dout[712]=40'b0;
dout[713]=40'b0;
dout[714]=40'b0;
dout[715]=40'b0;
dout[716]=40'b0;
dout[717]=40'b0;
dout[718]=40'b0;
dout[719]=40'b0;
dout[720]=40'b0;
dout[721]=40'b0;
dout[722]=40'b0;
dout[723]=40'b0;
dout[724]=40'b0;
dout[725]=40'b0;
dout[726]=40'b0;
dout[727]=40'b0;
dout[728]=40'b0;
dout[729]=40'b0;
dout[730]=40'b0;
dout[731]=40'b0;
dout[732]=40'b0;
dout[733]=40'b0;
dout[734]=40'b0;
dout[735]=40'b0;
dout[736]=40'b0;
dout[737]=40'b0;
dout[738]=40'b0;
dout[739]=40'b0;
dout[740]=40'b0;
dout[741]=40'b0;
dout[742]=40'b0;
dout[743]=40'b0;
dout[744]=40'b0;
dout[745]=40'b0;
dout[746]=40'b0;
dout[747]=40'b0;
dout[748]=40'b0;
dout[749]=40'b0;
dout[750]=40'b0;
dout[751]=40'b0;
dout[752]=40'b0;
dout[753]=40'b0;
dout[754]=40'b0;
dout[755]=40'b0;
dout[756]=40'b0;
dout[757]=40'b0;
dout[758]=40'b0;
dout[759]=40'b0;
dout[760]=40'b0;
dout[761]=40'b0;
dout[762]=40'b0;
dout[763]=40'b0;
dout[764]=40'b0;
dout[765]=40'b0;
dout[766]=40'b0;
dout[767]=40'b0;
dout[768]=40'b0;
dout[769]=40'b0;
dout[770]=40'b0;
dout[771]=40'b0;
dout[772]=40'b0;
dout[773]=40'b0;
dout[774]=40'b0;
dout[775]=40'b0;
dout[776]=40'b0;
dout[777]=40'b0;
dout[778]=40'b0;
dout[779]=40'b0;
dout[780]=40'b0;
dout[781]=40'b0;
dout[782]=40'b0;
dout[783]=40'b0;
dout[784]=40'b0;
dout[785]=40'b0;
dout[786]=40'b0;
dout[787]=40'b0;
dout[788]=40'b0;
dout[789]=40'b0;
dout[790]=40'b0;
dout[791]=40'b0;
dout[792]=40'b0;
dout[793]=40'b0;
dout[794]=40'b0;
dout[795]=40'b0;
dout[796]=40'b0;
dout[797]=40'b0;
dout[798]=40'b0;
dout[799]=40'b0;
dout[800]=40'b0;
dout[801]=40'b0;
dout[802]=40'b0;
dout[803]=40'b0;
dout[804]=40'b0;
dout[805]=40'b0;
dout[806]=40'b0;
dout[807]=40'b0;
dout[808]=40'b0;
dout[809]=40'b0;
dout[810]=40'b0;
dout[811]=40'b0;
dout[812]=40'b0;
dout[813]=40'b0;
dout[814]=40'b0;
dout[815]=40'b0;
dout[816]=40'b0;
dout[817]=40'b0;
dout[818]=40'b0;
dout[819]=40'b0;
dout[820]=40'b0;
dout[821]=40'b0;
dout[822]=40'b0;
dout[823]=40'b0;
dout[824]=40'b0;
dout[825]=40'b0;
dout[826]=40'b0;
dout[827]=40'b0;
dout[828]=40'b0;
dout[829]=40'b0;
dout[830]=40'b0;
dout[831]=40'b0;
dout[832]=40'b0;
dout[833]=40'b0;
dout[834]=40'b0;
dout[835]=40'b0;
dout[836]=40'b0;
dout[837]=40'b0;
dout[838]=40'b0;
dout[839]=40'b0;
dout[840]=40'b0;
dout[841]=40'b0;
dout[842]=40'b0;
dout[843]=40'b0;
dout[844]=40'b0;
dout[845]=40'b0;
dout[846]=40'b0;
dout[847]=40'b0;
dout[848]=40'b0;
dout[849]=40'b0;
dout[850]=40'b0;
dout[851]=40'b0;
dout[852]=40'b0;
dout[853]=40'b0;
dout[854]=40'b0;
dout[855]=40'b0;
dout[856]=40'b0;
dout[857]=40'b0;
dout[858]=40'b0;
dout[859]=40'b0;
dout[860]=40'b0;
dout[861]=40'b0;
dout[862]=40'b0;
dout[863]=40'b0;
dout[864]=40'b0;
dout[865]=40'b0;
dout[866]=40'b0;
dout[867]=40'b0;
dout[868]=40'b0;
dout[869]=40'b0;
dout[870]=40'b0;
dout[871]=40'b0;
dout[872]=40'b0;
dout[873]=40'b0;
dout[874]=40'b0;
dout[875]=40'b0;
dout[876]=40'b0;
dout[877]=40'b0;
dout[878]=40'b0;
dout[879]=40'b0;
dout[880]=40'b0;
dout[881]=40'b0;
dout[882]=40'b0;
dout[883]=40'b0;
dout[884]=40'b0;
dout[885]=40'b0;
dout[886]=40'b0;
dout[887]=40'b0;
dout[888]=40'b0;
dout[889]=40'b0;
dout[890]=40'b0;
dout[891]=40'b0;
dout[892]=40'b0;
dout[893]=40'b0;
dout[894]=40'b0;
dout[895]=40'b0;
dout[896]=40'b0;
dout[897]=40'b0;
dout[898]=40'b0;
dout[899]=40'b0;
dout[900]=40'b0;
dout[901]=40'b0;
dout[902]=40'b0;
dout[903]=40'b0;
dout[904]=40'b0;
dout[905]=40'b0;
dout[906]=40'b0;
dout[907]=40'b0;
dout[908]=40'b0;
dout[909]=40'b0;
dout[910]=40'b0;
dout[911]=40'b0;
dout[912]=40'b0;
dout[913]=40'b0;
dout[914]=40'b0;
dout[915]=40'b0;
dout[916]=40'b0;
dout[917]=40'b0;
dout[918]=40'b0;
dout[919]=40'b0;
dout[920]=40'b0;
dout[921]=40'b0;
dout[922]=40'b0;
dout[923]=40'b0;
dout[924]=40'b0;
dout[925]=40'b0;
dout[926]=40'b0;
dout[927]=40'b0;
dout[928]=40'b0;
dout[929]=40'b0;
dout[930]=40'b0;
dout[931]=40'b0;
dout[932]=40'b0;
dout[933]=40'b0;
dout[934]=40'b0;
dout[935]=40'b0;
dout[936]=40'b0;
dout[937]=40'b0;
dout[938]=40'b0;
dout[939]=40'b0;
dout[940]=40'b0;
dout[941]=40'b0;
dout[942]=40'b0;
dout[943]=40'b0;
dout[944]=40'b0;
dout[945]=40'b0;
dout[946]=40'b0;
dout[947]=40'b0;
dout[948]=40'b0;
dout[949]=40'b0;
dout[950]=40'b0;
dout[951]=40'b0;
dout[952]=40'b0;
dout[953]=40'b0;
dout[954]=40'b0;
dout[955]=40'b0;
dout[956]=40'b0;
dout[957]=40'b0;
dout[958]=40'b0;
dout[959]=40'b0;
dout[960]=40'b0;
dout[961]=40'b0;
dout[962]=40'b0;
dout[963]=40'b0;
dout[964]=40'b0;
dout[965]=40'b0;
dout[966]=40'b0;
dout[967]=40'b0;
dout[968]=40'b0;
dout[969]=40'b0;
dout[970]=40'b0;
dout[971]=40'b0;
dout[972]=40'b0;
dout[973]=40'b0;
dout[974]=40'b0;
dout[975]=40'b0;
dout[976]=40'b0;
dout[977]=40'b0;
dout[978]=40'b0;
dout[979]=40'b0;
dout[980]=40'b0;
dout[981]=40'b0;
dout[982]=40'b0;
dout[983]=40'b0;
dout[984]=40'b0;
dout[985]=40'b0;
dout[986]=40'b0;
dout[987]=40'b0;
dout[988]=40'b0;
dout[989]=40'b0;
dout[990]=40'b0;
dout[991]=40'b0;
dout[992]=40'b0;
dout[993]=40'b0;
dout[994]=40'b0;
dout[995]=40'b0;
dout[996]=40'b0;
dout[997]=40'b0;
dout[998]=40'b0;
dout[999]=40'b0;
dout[1000]=40'b0;
dout[1001]=40'b0;
dout[1002]=40'b0;
dout[1003]=40'b0;
dout[1004]=40'b0;
dout[1005]=40'b0;
dout[1006]=40'b0;
dout[1007]=40'b0;
dout[1008]=40'b0;
dout[1009]=40'b0;
dout[1010]=40'b0;
dout[1011]=40'b0;
dout[1012]=40'b0;
dout[1013]=40'b0;
dout[1014]=40'b0;
dout[1015]=40'b0;
dout[1016]=40'b0;
dout[1017]=40'b0;
dout[1018]=40'b0;
dout[1019]=40'b0;
dout[1020]=40'b0;
dout[1021]=40'b0;
dout[1022]=40'b0;
dout[1023]=40'b0;
end

always @ (posedge clk) begin
  w <= dout[addr];
end


endmodule

/** @} */ /* End of addtogroup ModMiscIpDspFftR22Sdc */
/* END OF FILE */